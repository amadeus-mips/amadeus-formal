module LUTRam(
  input         clock,
  input         reset,
  input  [7:0]  io_readAddr,
  output [20:0] io_readData,
  input  [7:0]  io_writeAddr,
  input  [20:0] io_writeData,
  input         io_writeEnable
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
`endif // RANDOMIZE_REG_INIT
  reg [20:0] _T_1_0; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_1; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_2; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_3; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_4; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_5; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_6; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_7; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_8; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_9; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_10; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_11; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_12; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_13; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_14; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_15; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_16; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_17; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_18; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_19; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_20; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_21; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_22; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_23; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_24; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_25; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_26; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_27; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_28; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_29; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_30; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_31; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_32; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_33; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_34; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_35; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_36; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_37; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_38; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_39; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_40; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_41; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_42; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_43; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_44; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_45; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_46; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_47; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_48; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_49; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_50; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_51; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_52; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_53; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_54; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_55; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_56; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_57; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_58; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_59; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_60; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_61; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_62; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_63; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_64; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_65; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_66; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_67; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_68; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_69; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_70; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_71; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_72; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_73; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_74; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_75; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_76; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_77; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_78; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_79; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_80; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_81; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_82; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_83; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_84; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_85; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_86; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_87; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_88; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_89; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_90; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_91; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_92; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_93; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_94; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_95; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_96; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_97; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_98; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_99; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_100; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_101; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_102; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_103; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_104; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_105; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_106; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_107; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_108; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_109; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_110; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_111; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_112; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_113; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_114; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_115; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_116; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_117; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_118; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_119; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_120; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_121; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_122; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_123; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_124; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_125; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_126; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_127; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_128; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_129; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_130; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_131; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_132; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_133; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_134; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_135; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_136; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_137; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_138; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_139; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_140; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_141; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_142; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_143; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_144; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_145; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_146; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_147; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_148; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_149; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_150; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_151; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_152; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_153; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_154; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_155; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_156; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_157; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_158; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_159; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_160; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_161; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_162; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_163; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_164; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_165; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_166; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_167; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_168; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_169; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_170; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_171; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_172; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_173; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_174; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_175; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_176; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_177; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_178; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_179; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_180; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_181; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_182; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_183; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_184; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_185; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_186; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_187; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_188; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_189; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_190; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_191; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_192; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_193; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_194; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_195; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_196; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_197; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_198; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_199; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_200; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_201; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_202; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_203; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_204; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_205; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_206; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_207; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_208; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_209; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_210; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_211; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_212; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_213; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_214; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_215; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_216; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_217; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_218; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_219; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_220; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_221; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_222; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_223; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_224; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_225; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_226; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_227; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_228; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_229; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_230; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_231; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_232; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_233; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_234; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_235; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_236; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_237; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_238; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_239; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_240; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_241; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_242; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_243; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_244; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_245; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_246; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_247; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_248; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_249; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_250; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_251; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_252; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_253; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_254; // @[LUTRam.scala 57:19]
  reg [20:0] _T_1_255; // @[LUTRam.scala 57:19]
  wire [20:0] _GEN_1 = 8'h1 == io_readAddr ? _T_1_1 : _T_1_0; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_2 = 8'h2 == io_readAddr ? _T_1_2 : _GEN_1; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_3 = 8'h3 == io_readAddr ? _T_1_3 : _GEN_2; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_4 = 8'h4 == io_readAddr ? _T_1_4 : _GEN_3; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_5 = 8'h5 == io_readAddr ? _T_1_5 : _GEN_4; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_6 = 8'h6 == io_readAddr ? _T_1_6 : _GEN_5; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_7 = 8'h7 == io_readAddr ? _T_1_7 : _GEN_6; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_8 = 8'h8 == io_readAddr ? _T_1_8 : _GEN_7; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_9 = 8'h9 == io_readAddr ? _T_1_9 : _GEN_8; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_10 = 8'ha == io_readAddr ? _T_1_10 : _GEN_9; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_11 = 8'hb == io_readAddr ? _T_1_11 : _GEN_10; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_12 = 8'hc == io_readAddr ? _T_1_12 : _GEN_11; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_13 = 8'hd == io_readAddr ? _T_1_13 : _GEN_12; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_14 = 8'he == io_readAddr ? _T_1_14 : _GEN_13; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_15 = 8'hf == io_readAddr ? _T_1_15 : _GEN_14; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_16 = 8'h10 == io_readAddr ? _T_1_16 : _GEN_15; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_17 = 8'h11 == io_readAddr ? _T_1_17 : _GEN_16; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_18 = 8'h12 == io_readAddr ? _T_1_18 : _GEN_17; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_19 = 8'h13 == io_readAddr ? _T_1_19 : _GEN_18; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_20 = 8'h14 == io_readAddr ? _T_1_20 : _GEN_19; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_21 = 8'h15 == io_readAddr ? _T_1_21 : _GEN_20; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_22 = 8'h16 == io_readAddr ? _T_1_22 : _GEN_21; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_23 = 8'h17 == io_readAddr ? _T_1_23 : _GEN_22; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_24 = 8'h18 == io_readAddr ? _T_1_24 : _GEN_23; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_25 = 8'h19 == io_readAddr ? _T_1_25 : _GEN_24; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_26 = 8'h1a == io_readAddr ? _T_1_26 : _GEN_25; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_27 = 8'h1b == io_readAddr ? _T_1_27 : _GEN_26; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_28 = 8'h1c == io_readAddr ? _T_1_28 : _GEN_27; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_29 = 8'h1d == io_readAddr ? _T_1_29 : _GEN_28; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_30 = 8'h1e == io_readAddr ? _T_1_30 : _GEN_29; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_31 = 8'h1f == io_readAddr ? _T_1_31 : _GEN_30; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_32 = 8'h20 == io_readAddr ? _T_1_32 : _GEN_31; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_33 = 8'h21 == io_readAddr ? _T_1_33 : _GEN_32; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_34 = 8'h22 == io_readAddr ? _T_1_34 : _GEN_33; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_35 = 8'h23 == io_readAddr ? _T_1_35 : _GEN_34; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_36 = 8'h24 == io_readAddr ? _T_1_36 : _GEN_35; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_37 = 8'h25 == io_readAddr ? _T_1_37 : _GEN_36; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_38 = 8'h26 == io_readAddr ? _T_1_38 : _GEN_37; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_39 = 8'h27 == io_readAddr ? _T_1_39 : _GEN_38; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_40 = 8'h28 == io_readAddr ? _T_1_40 : _GEN_39; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_41 = 8'h29 == io_readAddr ? _T_1_41 : _GEN_40; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_42 = 8'h2a == io_readAddr ? _T_1_42 : _GEN_41; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_43 = 8'h2b == io_readAddr ? _T_1_43 : _GEN_42; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_44 = 8'h2c == io_readAddr ? _T_1_44 : _GEN_43; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_45 = 8'h2d == io_readAddr ? _T_1_45 : _GEN_44; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_46 = 8'h2e == io_readAddr ? _T_1_46 : _GEN_45; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_47 = 8'h2f == io_readAddr ? _T_1_47 : _GEN_46; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_48 = 8'h30 == io_readAddr ? _T_1_48 : _GEN_47; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_49 = 8'h31 == io_readAddr ? _T_1_49 : _GEN_48; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_50 = 8'h32 == io_readAddr ? _T_1_50 : _GEN_49; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_51 = 8'h33 == io_readAddr ? _T_1_51 : _GEN_50; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_52 = 8'h34 == io_readAddr ? _T_1_52 : _GEN_51; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_53 = 8'h35 == io_readAddr ? _T_1_53 : _GEN_52; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_54 = 8'h36 == io_readAddr ? _T_1_54 : _GEN_53; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_55 = 8'h37 == io_readAddr ? _T_1_55 : _GEN_54; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_56 = 8'h38 == io_readAddr ? _T_1_56 : _GEN_55; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_57 = 8'h39 == io_readAddr ? _T_1_57 : _GEN_56; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_58 = 8'h3a == io_readAddr ? _T_1_58 : _GEN_57; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_59 = 8'h3b == io_readAddr ? _T_1_59 : _GEN_58; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_60 = 8'h3c == io_readAddr ? _T_1_60 : _GEN_59; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_61 = 8'h3d == io_readAddr ? _T_1_61 : _GEN_60; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_62 = 8'h3e == io_readAddr ? _T_1_62 : _GEN_61; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_63 = 8'h3f == io_readAddr ? _T_1_63 : _GEN_62; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_64 = 8'h40 == io_readAddr ? _T_1_64 : _GEN_63; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_65 = 8'h41 == io_readAddr ? _T_1_65 : _GEN_64; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_66 = 8'h42 == io_readAddr ? _T_1_66 : _GEN_65; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_67 = 8'h43 == io_readAddr ? _T_1_67 : _GEN_66; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_68 = 8'h44 == io_readAddr ? _T_1_68 : _GEN_67; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_69 = 8'h45 == io_readAddr ? _T_1_69 : _GEN_68; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_70 = 8'h46 == io_readAddr ? _T_1_70 : _GEN_69; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_71 = 8'h47 == io_readAddr ? _T_1_71 : _GEN_70; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_72 = 8'h48 == io_readAddr ? _T_1_72 : _GEN_71; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_73 = 8'h49 == io_readAddr ? _T_1_73 : _GEN_72; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_74 = 8'h4a == io_readAddr ? _T_1_74 : _GEN_73; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_75 = 8'h4b == io_readAddr ? _T_1_75 : _GEN_74; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_76 = 8'h4c == io_readAddr ? _T_1_76 : _GEN_75; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_77 = 8'h4d == io_readAddr ? _T_1_77 : _GEN_76; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_78 = 8'h4e == io_readAddr ? _T_1_78 : _GEN_77; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_79 = 8'h4f == io_readAddr ? _T_1_79 : _GEN_78; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_80 = 8'h50 == io_readAddr ? _T_1_80 : _GEN_79; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_81 = 8'h51 == io_readAddr ? _T_1_81 : _GEN_80; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_82 = 8'h52 == io_readAddr ? _T_1_82 : _GEN_81; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_83 = 8'h53 == io_readAddr ? _T_1_83 : _GEN_82; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_84 = 8'h54 == io_readAddr ? _T_1_84 : _GEN_83; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_85 = 8'h55 == io_readAddr ? _T_1_85 : _GEN_84; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_86 = 8'h56 == io_readAddr ? _T_1_86 : _GEN_85; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_87 = 8'h57 == io_readAddr ? _T_1_87 : _GEN_86; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_88 = 8'h58 == io_readAddr ? _T_1_88 : _GEN_87; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_89 = 8'h59 == io_readAddr ? _T_1_89 : _GEN_88; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_90 = 8'h5a == io_readAddr ? _T_1_90 : _GEN_89; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_91 = 8'h5b == io_readAddr ? _T_1_91 : _GEN_90; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_92 = 8'h5c == io_readAddr ? _T_1_92 : _GEN_91; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_93 = 8'h5d == io_readAddr ? _T_1_93 : _GEN_92; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_94 = 8'h5e == io_readAddr ? _T_1_94 : _GEN_93; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_95 = 8'h5f == io_readAddr ? _T_1_95 : _GEN_94; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_96 = 8'h60 == io_readAddr ? _T_1_96 : _GEN_95; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_97 = 8'h61 == io_readAddr ? _T_1_97 : _GEN_96; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_98 = 8'h62 == io_readAddr ? _T_1_98 : _GEN_97; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_99 = 8'h63 == io_readAddr ? _T_1_99 : _GEN_98; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_100 = 8'h64 == io_readAddr ? _T_1_100 : _GEN_99; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_101 = 8'h65 == io_readAddr ? _T_1_101 : _GEN_100; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_102 = 8'h66 == io_readAddr ? _T_1_102 : _GEN_101; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_103 = 8'h67 == io_readAddr ? _T_1_103 : _GEN_102; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_104 = 8'h68 == io_readAddr ? _T_1_104 : _GEN_103; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_105 = 8'h69 == io_readAddr ? _T_1_105 : _GEN_104; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_106 = 8'h6a == io_readAddr ? _T_1_106 : _GEN_105; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_107 = 8'h6b == io_readAddr ? _T_1_107 : _GEN_106; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_108 = 8'h6c == io_readAddr ? _T_1_108 : _GEN_107; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_109 = 8'h6d == io_readAddr ? _T_1_109 : _GEN_108; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_110 = 8'h6e == io_readAddr ? _T_1_110 : _GEN_109; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_111 = 8'h6f == io_readAddr ? _T_1_111 : _GEN_110; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_112 = 8'h70 == io_readAddr ? _T_1_112 : _GEN_111; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_113 = 8'h71 == io_readAddr ? _T_1_113 : _GEN_112; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_114 = 8'h72 == io_readAddr ? _T_1_114 : _GEN_113; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_115 = 8'h73 == io_readAddr ? _T_1_115 : _GEN_114; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_116 = 8'h74 == io_readAddr ? _T_1_116 : _GEN_115; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_117 = 8'h75 == io_readAddr ? _T_1_117 : _GEN_116; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_118 = 8'h76 == io_readAddr ? _T_1_118 : _GEN_117; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_119 = 8'h77 == io_readAddr ? _T_1_119 : _GEN_118; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_120 = 8'h78 == io_readAddr ? _T_1_120 : _GEN_119; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_121 = 8'h79 == io_readAddr ? _T_1_121 : _GEN_120; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_122 = 8'h7a == io_readAddr ? _T_1_122 : _GEN_121; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_123 = 8'h7b == io_readAddr ? _T_1_123 : _GEN_122; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_124 = 8'h7c == io_readAddr ? _T_1_124 : _GEN_123; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_125 = 8'h7d == io_readAddr ? _T_1_125 : _GEN_124; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_126 = 8'h7e == io_readAddr ? _T_1_126 : _GEN_125; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_127 = 8'h7f == io_readAddr ? _T_1_127 : _GEN_126; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_128 = 8'h80 == io_readAddr ? _T_1_128 : _GEN_127; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_129 = 8'h81 == io_readAddr ? _T_1_129 : _GEN_128; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_130 = 8'h82 == io_readAddr ? _T_1_130 : _GEN_129; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_131 = 8'h83 == io_readAddr ? _T_1_131 : _GEN_130; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_132 = 8'h84 == io_readAddr ? _T_1_132 : _GEN_131; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_133 = 8'h85 == io_readAddr ? _T_1_133 : _GEN_132; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_134 = 8'h86 == io_readAddr ? _T_1_134 : _GEN_133; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_135 = 8'h87 == io_readAddr ? _T_1_135 : _GEN_134; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_136 = 8'h88 == io_readAddr ? _T_1_136 : _GEN_135; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_137 = 8'h89 == io_readAddr ? _T_1_137 : _GEN_136; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_138 = 8'h8a == io_readAddr ? _T_1_138 : _GEN_137; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_139 = 8'h8b == io_readAddr ? _T_1_139 : _GEN_138; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_140 = 8'h8c == io_readAddr ? _T_1_140 : _GEN_139; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_141 = 8'h8d == io_readAddr ? _T_1_141 : _GEN_140; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_142 = 8'h8e == io_readAddr ? _T_1_142 : _GEN_141; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_143 = 8'h8f == io_readAddr ? _T_1_143 : _GEN_142; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_144 = 8'h90 == io_readAddr ? _T_1_144 : _GEN_143; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_145 = 8'h91 == io_readAddr ? _T_1_145 : _GEN_144; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_146 = 8'h92 == io_readAddr ? _T_1_146 : _GEN_145; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_147 = 8'h93 == io_readAddr ? _T_1_147 : _GEN_146; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_148 = 8'h94 == io_readAddr ? _T_1_148 : _GEN_147; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_149 = 8'h95 == io_readAddr ? _T_1_149 : _GEN_148; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_150 = 8'h96 == io_readAddr ? _T_1_150 : _GEN_149; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_151 = 8'h97 == io_readAddr ? _T_1_151 : _GEN_150; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_152 = 8'h98 == io_readAddr ? _T_1_152 : _GEN_151; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_153 = 8'h99 == io_readAddr ? _T_1_153 : _GEN_152; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_154 = 8'h9a == io_readAddr ? _T_1_154 : _GEN_153; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_155 = 8'h9b == io_readAddr ? _T_1_155 : _GEN_154; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_156 = 8'h9c == io_readAddr ? _T_1_156 : _GEN_155; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_157 = 8'h9d == io_readAddr ? _T_1_157 : _GEN_156; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_158 = 8'h9e == io_readAddr ? _T_1_158 : _GEN_157; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_159 = 8'h9f == io_readAddr ? _T_1_159 : _GEN_158; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_160 = 8'ha0 == io_readAddr ? _T_1_160 : _GEN_159; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_161 = 8'ha1 == io_readAddr ? _T_1_161 : _GEN_160; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_162 = 8'ha2 == io_readAddr ? _T_1_162 : _GEN_161; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_163 = 8'ha3 == io_readAddr ? _T_1_163 : _GEN_162; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_164 = 8'ha4 == io_readAddr ? _T_1_164 : _GEN_163; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_165 = 8'ha5 == io_readAddr ? _T_1_165 : _GEN_164; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_166 = 8'ha6 == io_readAddr ? _T_1_166 : _GEN_165; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_167 = 8'ha7 == io_readAddr ? _T_1_167 : _GEN_166; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_168 = 8'ha8 == io_readAddr ? _T_1_168 : _GEN_167; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_169 = 8'ha9 == io_readAddr ? _T_1_169 : _GEN_168; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_170 = 8'haa == io_readAddr ? _T_1_170 : _GEN_169; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_171 = 8'hab == io_readAddr ? _T_1_171 : _GEN_170; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_172 = 8'hac == io_readAddr ? _T_1_172 : _GEN_171; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_173 = 8'had == io_readAddr ? _T_1_173 : _GEN_172; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_174 = 8'hae == io_readAddr ? _T_1_174 : _GEN_173; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_175 = 8'haf == io_readAddr ? _T_1_175 : _GEN_174; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_176 = 8'hb0 == io_readAddr ? _T_1_176 : _GEN_175; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_177 = 8'hb1 == io_readAddr ? _T_1_177 : _GEN_176; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_178 = 8'hb2 == io_readAddr ? _T_1_178 : _GEN_177; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_179 = 8'hb3 == io_readAddr ? _T_1_179 : _GEN_178; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_180 = 8'hb4 == io_readAddr ? _T_1_180 : _GEN_179; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_181 = 8'hb5 == io_readAddr ? _T_1_181 : _GEN_180; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_182 = 8'hb6 == io_readAddr ? _T_1_182 : _GEN_181; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_183 = 8'hb7 == io_readAddr ? _T_1_183 : _GEN_182; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_184 = 8'hb8 == io_readAddr ? _T_1_184 : _GEN_183; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_185 = 8'hb9 == io_readAddr ? _T_1_185 : _GEN_184; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_186 = 8'hba == io_readAddr ? _T_1_186 : _GEN_185; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_187 = 8'hbb == io_readAddr ? _T_1_187 : _GEN_186; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_188 = 8'hbc == io_readAddr ? _T_1_188 : _GEN_187; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_189 = 8'hbd == io_readAddr ? _T_1_189 : _GEN_188; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_190 = 8'hbe == io_readAddr ? _T_1_190 : _GEN_189; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_191 = 8'hbf == io_readAddr ? _T_1_191 : _GEN_190; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_192 = 8'hc0 == io_readAddr ? _T_1_192 : _GEN_191; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_193 = 8'hc1 == io_readAddr ? _T_1_193 : _GEN_192; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_194 = 8'hc2 == io_readAddr ? _T_1_194 : _GEN_193; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_195 = 8'hc3 == io_readAddr ? _T_1_195 : _GEN_194; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_196 = 8'hc4 == io_readAddr ? _T_1_196 : _GEN_195; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_197 = 8'hc5 == io_readAddr ? _T_1_197 : _GEN_196; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_198 = 8'hc6 == io_readAddr ? _T_1_198 : _GEN_197; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_199 = 8'hc7 == io_readAddr ? _T_1_199 : _GEN_198; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_200 = 8'hc8 == io_readAddr ? _T_1_200 : _GEN_199; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_201 = 8'hc9 == io_readAddr ? _T_1_201 : _GEN_200; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_202 = 8'hca == io_readAddr ? _T_1_202 : _GEN_201; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_203 = 8'hcb == io_readAddr ? _T_1_203 : _GEN_202; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_204 = 8'hcc == io_readAddr ? _T_1_204 : _GEN_203; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_205 = 8'hcd == io_readAddr ? _T_1_205 : _GEN_204; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_206 = 8'hce == io_readAddr ? _T_1_206 : _GEN_205; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_207 = 8'hcf == io_readAddr ? _T_1_207 : _GEN_206; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_208 = 8'hd0 == io_readAddr ? _T_1_208 : _GEN_207; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_209 = 8'hd1 == io_readAddr ? _T_1_209 : _GEN_208; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_210 = 8'hd2 == io_readAddr ? _T_1_210 : _GEN_209; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_211 = 8'hd3 == io_readAddr ? _T_1_211 : _GEN_210; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_212 = 8'hd4 == io_readAddr ? _T_1_212 : _GEN_211; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_213 = 8'hd5 == io_readAddr ? _T_1_213 : _GEN_212; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_214 = 8'hd6 == io_readAddr ? _T_1_214 : _GEN_213; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_215 = 8'hd7 == io_readAddr ? _T_1_215 : _GEN_214; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_216 = 8'hd8 == io_readAddr ? _T_1_216 : _GEN_215; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_217 = 8'hd9 == io_readAddr ? _T_1_217 : _GEN_216; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_218 = 8'hda == io_readAddr ? _T_1_218 : _GEN_217; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_219 = 8'hdb == io_readAddr ? _T_1_219 : _GEN_218; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_220 = 8'hdc == io_readAddr ? _T_1_220 : _GEN_219; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_221 = 8'hdd == io_readAddr ? _T_1_221 : _GEN_220; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_222 = 8'hde == io_readAddr ? _T_1_222 : _GEN_221; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_223 = 8'hdf == io_readAddr ? _T_1_223 : _GEN_222; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_224 = 8'he0 == io_readAddr ? _T_1_224 : _GEN_223; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_225 = 8'he1 == io_readAddr ? _T_1_225 : _GEN_224; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_226 = 8'he2 == io_readAddr ? _T_1_226 : _GEN_225; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_227 = 8'he3 == io_readAddr ? _T_1_227 : _GEN_226; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_228 = 8'he4 == io_readAddr ? _T_1_228 : _GEN_227; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_229 = 8'he5 == io_readAddr ? _T_1_229 : _GEN_228; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_230 = 8'he6 == io_readAddr ? _T_1_230 : _GEN_229; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_231 = 8'he7 == io_readAddr ? _T_1_231 : _GEN_230; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_232 = 8'he8 == io_readAddr ? _T_1_232 : _GEN_231; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_233 = 8'he9 == io_readAddr ? _T_1_233 : _GEN_232; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_234 = 8'hea == io_readAddr ? _T_1_234 : _GEN_233; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_235 = 8'heb == io_readAddr ? _T_1_235 : _GEN_234; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_236 = 8'hec == io_readAddr ? _T_1_236 : _GEN_235; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_237 = 8'hed == io_readAddr ? _T_1_237 : _GEN_236; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_238 = 8'hee == io_readAddr ? _T_1_238 : _GEN_237; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_239 = 8'hef == io_readAddr ? _T_1_239 : _GEN_238; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_240 = 8'hf0 == io_readAddr ? _T_1_240 : _GEN_239; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_241 = 8'hf1 == io_readAddr ? _T_1_241 : _GEN_240; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_242 = 8'hf2 == io_readAddr ? _T_1_242 : _GEN_241; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_243 = 8'hf3 == io_readAddr ? _T_1_243 : _GEN_242; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_244 = 8'hf4 == io_readAddr ? _T_1_244 : _GEN_243; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_245 = 8'hf5 == io_readAddr ? _T_1_245 : _GEN_244; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_246 = 8'hf6 == io_readAddr ? _T_1_246 : _GEN_245; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_247 = 8'hf7 == io_readAddr ? _T_1_247 : _GEN_246; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_248 = 8'hf8 == io_readAddr ? _T_1_248 : _GEN_247; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_249 = 8'hf9 == io_readAddr ? _T_1_249 : _GEN_248; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_250 = 8'hfa == io_readAddr ? _T_1_250 : _GEN_249; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_251 = 8'hfb == io_readAddr ? _T_1_251 : _GEN_250; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_252 = 8'hfc == io_readAddr ? _T_1_252 : _GEN_251; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_253 = 8'hfd == io_readAddr ? _T_1_253 : _GEN_252; // @[LUTRam.scala 58:20]
  wire [20:0] _GEN_254 = 8'hfe == io_readAddr ? _T_1_254 : _GEN_253; // @[LUTRam.scala 58:20]
  assign io_readData = 8'hff == io_readAddr ? _T_1_255 : _GEN_254; // @[LUTRam.scala 58:20]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_1_0 = _RAND_0[20:0];
  _RAND_1 = {1{`RANDOM}};
  _T_1_1 = _RAND_1[20:0];
  _RAND_2 = {1{`RANDOM}};
  _T_1_2 = _RAND_2[20:0];
  _RAND_3 = {1{`RANDOM}};
  _T_1_3 = _RAND_3[20:0];
  _RAND_4 = {1{`RANDOM}};
  _T_1_4 = _RAND_4[20:0];
  _RAND_5 = {1{`RANDOM}};
  _T_1_5 = _RAND_5[20:0];
  _RAND_6 = {1{`RANDOM}};
  _T_1_6 = _RAND_6[20:0];
  _RAND_7 = {1{`RANDOM}};
  _T_1_7 = _RAND_7[20:0];
  _RAND_8 = {1{`RANDOM}};
  _T_1_8 = _RAND_8[20:0];
  _RAND_9 = {1{`RANDOM}};
  _T_1_9 = _RAND_9[20:0];
  _RAND_10 = {1{`RANDOM}};
  _T_1_10 = _RAND_10[20:0];
  _RAND_11 = {1{`RANDOM}};
  _T_1_11 = _RAND_11[20:0];
  _RAND_12 = {1{`RANDOM}};
  _T_1_12 = _RAND_12[20:0];
  _RAND_13 = {1{`RANDOM}};
  _T_1_13 = _RAND_13[20:0];
  _RAND_14 = {1{`RANDOM}};
  _T_1_14 = _RAND_14[20:0];
  _RAND_15 = {1{`RANDOM}};
  _T_1_15 = _RAND_15[20:0];
  _RAND_16 = {1{`RANDOM}};
  _T_1_16 = _RAND_16[20:0];
  _RAND_17 = {1{`RANDOM}};
  _T_1_17 = _RAND_17[20:0];
  _RAND_18 = {1{`RANDOM}};
  _T_1_18 = _RAND_18[20:0];
  _RAND_19 = {1{`RANDOM}};
  _T_1_19 = _RAND_19[20:0];
  _RAND_20 = {1{`RANDOM}};
  _T_1_20 = _RAND_20[20:0];
  _RAND_21 = {1{`RANDOM}};
  _T_1_21 = _RAND_21[20:0];
  _RAND_22 = {1{`RANDOM}};
  _T_1_22 = _RAND_22[20:0];
  _RAND_23 = {1{`RANDOM}};
  _T_1_23 = _RAND_23[20:0];
  _RAND_24 = {1{`RANDOM}};
  _T_1_24 = _RAND_24[20:0];
  _RAND_25 = {1{`RANDOM}};
  _T_1_25 = _RAND_25[20:0];
  _RAND_26 = {1{`RANDOM}};
  _T_1_26 = _RAND_26[20:0];
  _RAND_27 = {1{`RANDOM}};
  _T_1_27 = _RAND_27[20:0];
  _RAND_28 = {1{`RANDOM}};
  _T_1_28 = _RAND_28[20:0];
  _RAND_29 = {1{`RANDOM}};
  _T_1_29 = _RAND_29[20:0];
  _RAND_30 = {1{`RANDOM}};
  _T_1_30 = _RAND_30[20:0];
  _RAND_31 = {1{`RANDOM}};
  _T_1_31 = _RAND_31[20:0];
  _RAND_32 = {1{`RANDOM}};
  _T_1_32 = _RAND_32[20:0];
  _RAND_33 = {1{`RANDOM}};
  _T_1_33 = _RAND_33[20:0];
  _RAND_34 = {1{`RANDOM}};
  _T_1_34 = _RAND_34[20:0];
  _RAND_35 = {1{`RANDOM}};
  _T_1_35 = _RAND_35[20:0];
  _RAND_36 = {1{`RANDOM}};
  _T_1_36 = _RAND_36[20:0];
  _RAND_37 = {1{`RANDOM}};
  _T_1_37 = _RAND_37[20:0];
  _RAND_38 = {1{`RANDOM}};
  _T_1_38 = _RAND_38[20:0];
  _RAND_39 = {1{`RANDOM}};
  _T_1_39 = _RAND_39[20:0];
  _RAND_40 = {1{`RANDOM}};
  _T_1_40 = _RAND_40[20:0];
  _RAND_41 = {1{`RANDOM}};
  _T_1_41 = _RAND_41[20:0];
  _RAND_42 = {1{`RANDOM}};
  _T_1_42 = _RAND_42[20:0];
  _RAND_43 = {1{`RANDOM}};
  _T_1_43 = _RAND_43[20:0];
  _RAND_44 = {1{`RANDOM}};
  _T_1_44 = _RAND_44[20:0];
  _RAND_45 = {1{`RANDOM}};
  _T_1_45 = _RAND_45[20:0];
  _RAND_46 = {1{`RANDOM}};
  _T_1_46 = _RAND_46[20:0];
  _RAND_47 = {1{`RANDOM}};
  _T_1_47 = _RAND_47[20:0];
  _RAND_48 = {1{`RANDOM}};
  _T_1_48 = _RAND_48[20:0];
  _RAND_49 = {1{`RANDOM}};
  _T_1_49 = _RAND_49[20:0];
  _RAND_50 = {1{`RANDOM}};
  _T_1_50 = _RAND_50[20:0];
  _RAND_51 = {1{`RANDOM}};
  _T_1_51 = _RAND_51[20:0];
  _RAND_52 = {1{`RANDOM}};
  _T_1_52 = _RAND_52[20:0];
  _RAND_53 = {1{`RANDOM}};
  _T_1_53 = _RAND_53[20:0];
  _RAND_54 = {1{`RANDOM}};
  _T_1_54 = _RAND_54[20:0];
  _RAND_55 = {1{`RANDOM}};
  _T_1_55 = _RAND_55[20:0];
  _RAND_56 = {1{`RANDOM}};
  _T_1_56 = _RAND_56[20:0];
  _RAND_57 = {1{`RANDOM}};
  _T_1_57 = _RAND_57[20:0];
  _RAND_58 = {1{`RANDOM}};
  _T_1_58 = _RAND_58[20:0];
  _RAND_59 = {1{`RANDOM}};
  _T_1_59 = _RAND_59[20:0];
  _RAND_60 = {1{`RANDOM}};
  _T_1_60 = _RAND_60[20:0];
  _RAND_61 = {1{`RANDOM}};
  _T_1_61 = _RAND_61[20:0];
  _RAND_62 = {1{`RANDOM}};
  _T_1_62 = _RAND_62[20:0];
  _RAND_63 = {1{`RANDOM}};
  _T_1_63 = _RAND_63[20:0];
  _RAND_64 = {1{`RANDOM}};
  _T_1_64 = _RAND_64[20:0];
  _RAND_65 = {1{`RANDOM}};
  _T_1_65 = _RAND_65[20:0];
  _RAND_66 = {1{`RANDOM}};
  _T_1_66 = _RAND_66[20:0];
  _RAND_67 = {1{`RANDOM}};
  _T_1_67 = _RAND_67[20:0];
  _RAND_68 = {1{`RANDOM}};
  _T_1_68 = _RAND_68[20:0];
  _RAND_69 = {1{`RANDOM}};
  _T_1_69 = _RAND_69[20:0];
  _RAND_70 = {1{`RANDOM}};
  _T_1_70 = _RAND_70[20:0];
  _RAND_71 = {1{`RANDOM}};
  _T_1_71 = _RAND_71[20:0];
  _RAND_72 = {1{`RANDOM}};
  _T_1_72 = _RAND_72[20:0];
  _RAND_73 = {1{`RANDOM}};
  _T_1_73 = _RAND_73[20:0];
  _RAND_74 = {1{`RANDOM}};
  _T_1_74 = _RAND_74[20:0];
  _RAND_75 = {1{`RANDOM}};
  _T_1_75 = _RAND_75[20:0];
  _RAND_76 = {1{`RANDOM}};
  _T_1_76 = _RAND_76[20:0];
  _RAND_77 = {1{`RANDOM}};
  _T_1_77 = _RAND_77[20:0];
  _RAND_78 = {1{`RANDOM}};
  _T_1_78 = _RAND_78[20:0];
  _RAND_79 = {1{`RANDOM}};
  _T_1_79 = _RAND_79[20:0];
  _RAND_80 = {1{`RANDOM}};
  _T_1_80 = _RAND_80[20:0];
  _RAND_81 = {1{`RANDOM}};
  _T_1_81 = _RAND_81[20:0];
  _RAND_82 = {1{`RANDOM}};
  _T_1_82 = _RAND_82[20:0];
  _RAND_83 = {1{`RANDOM}};
  _T_1_83 = _RAND_83[20:0];
  _RAND_84 = {1{`RANDOM}};
  _T_1_84 = _RAND_84[20:0];
  _RAND_85 = {1{`RANDOM}};
  _T_1_85 = _RAND_85[20:0];
  _RAND_86 = {1{`RANDOM}};
  _T_1_86 = _RAND_86[20:0];
  _RAND_87 = {1{`RANDOM}};
  _T_1_87 = _RAND_87[20:0];
  _RAND_88 = {1{`RANDOM}};
  _T_1_88 = _RAND_88[20:0];
  _RAND_89 = {1{`RANDOM}};
  _T_1_89 = _RAND_89[20:0];
  _RAND_90 = {1{`RANDOM}};
  _T_1_90 = _RAND_90[20:0];
  _RAND_91 = {1{`RANDOM}};
  _T_1_91 = _RAND_91[20:0];
  _RAND_92 = {1{`RANDOM}};
  _T_1_92 = _RAND_92[20:0];
  _RAND_93 = {1{`RANDOM}};
  _T_1_93 = _RAND_93[20:0];
  _RAND_94 = {1{`RANDOM}};
  _T_1_94 = _RAND_94[20:0];
  _RAND_95 = {1{`RANDOM}};
  _T_1_95 = _RAND_95[20:0];
  _RAND_96 = {1{`RANDOM}};
  _T_1_96 = _RAND_96[20:0];
  _RAND_97 = {1{`RANDOM}};
  _T_1_97 = _RAND_97[20:0];
  _RAND_98 = {1{`RANDOM}};
  _T_1_98 = _RAND_98[20:0];
  _RAND_99 = {1{`RANDOM}};
  _T_1_99 = _RAND_99[20:0];
  _RAND_100 = {1{`RANDOM}};
  _T_1_100 = _RAND_100[20:0];
  _RAND_101 = {1{`RANDOM}};
  _T_1_101 = _RAND_101[20:0];
  _RAND_102 = {1{`RANDOM}};
  _T_1_102 = _RAND_102[20:0];
  _RAND_103 = {1{`RANDOM}};
  _T_1_103 = _RAND_103[20:0];
  _RAND_104 = {1{`RANDOM}};
  _T_1_104 = _RAND_104[20:0];
  _RAND_105 = {1{`RANDOM}};
  _T_1_105 = _RAND_105[20:0];
  _RAND_106 = {1{`RANDOM}};
  _T_1_106 = _RAND_106[20:0];
  _RAND_107 = {1{`RANDOM}};
  _T_1_107 = _RAND_107[20:0];
  _RAND_108 = {1{`RANDOM}};
  _T_1_108 = _RAND_108[20:0];
  _RAND_109 = {1{`RANDOM}};
  _T_1_109 = _RAND_109[20:0];
  _RAND_110 = {1{`RANDOM}};
  _T_1_110 = _RAND_110[20:0];
  _RAND_111 = {1{`RANDOM}};
  _T_1_111 = _RAND_111[20:0];
  _RAND_112 = {1{`RANDOM}};
  _T_1_112 = _RAND_112[20:0];
  _RAND_113 = {1{`RANDOM}};
  _T_1_113 = _RAND_113[20:0];
  _RAND_114 = {1{`RANDOM}};
  _T_1_114 = _RAND_114[20:0];
  _RAND_115 = {1{`RANDOM}};
  _T_1_115 = _RAND_115[20:0];
  _RAND_116 = {1{`RANDOM}};
  _T_1_116 = _RAND_116[20:0];
  _RAND_117 = {1{`RANDOM}};
  _T_1_117 = _RAND_117[20:0];
  _RAND_118 = {1{`RANDOM}};
  _T_1_118 = _RAND_118[20:0];
  _RAND_119 = {1{`RANDOM}};
  _T_1_119 = _RAND_119[20:0];
  _RAND_120 = {1{`RANDOM}};
  _T_1_120 = _RAND_120[20:0];
  _RAND_121 = {1{`RANDOM}};
  _T_1_121 = _RAND_121[20:0];
  _RAND_122 = {1{`RANDOM}};
  _T_1_122 = _RAND_122[20:0];
  _RAND_123 = {1{`RANDOM}};
  _T_1_123 = _RAND_123[20:0];
  _RAND_124 = {1{`RANDOM}};
  _T_1_124 = _RAND_124[20:0];
  _RAND_125 = {1{`RANDOM}};
  _T_1_125 = _RAND_125[20:0];
  _RAND_126 = {1{`RANDOM}};
  _T_1_126 = _RAND_126[20:0];
  _RAND_127 = {1{`RANDOM}};
  _T_1_127 = _RAND_127[20:0];
  _RAND_128 = {1{`RANDOM}};
  _T_1_128 = _RAND_128[20:0];
  _RAND_129 = {1{`RANDOM}};
  _T_1_129 = _RAND_129[20:0];
  _RAND_130 = {1{`RANDOM}};
  _T_1_130 = _RAND_130[20:0];
  _RAND_131 = {1{`RANDOM}};
  _T_1_131 = _RAND_131[20:0];
  _RAND_132 = {1{`RANDOM}};
  _T_1_132 = _RAND_132[20:0];
  _RAND_133 = {1{`RANDOM}};
  _T_1_133 = _RAND_133[20:0];
  _RAND_134 = {1{`RANDOM}};
  _T_1_134 = _RAND_134[20:0];
  _RAND_135 = {1{`RANDOM}};
  _T_1_135 = _RAND_135[20:0];
  _RAND_136 = {1{`RANDOM}};
  _T_1_136 = _RAND_136[20:0];
  _RAND_137 = {1{`RANDOM}};
  _T_1_137 = _RAND_137[20:0];
  _RAND_138 = {1{`RANDOM}};
  _T_1_138 = _RAND_138[20:0];
  _RAND_139 = {1{`RANDOM}};
  _T_1_139 = _RAND_139[20:0];
  _RAND_140 = {1{`RANDOM}};
  _T_1_140 = _RAND_140[20:0];
  _RAND_141 = {1{`RANDOM}};
  _T_1_141 = _RAND_141[20:0];
  _RAND_142 = {1{`RANDOM}};
  _T_1_142 = _RAND_142[20:0];
  _RAND_143 = {1{`RANDOM}};
  _T_1_143 = _RAND_143[20:0];
  _RAND_144 = {1{`RANDOM}};
  _T_1_144 = _RAND_144[20:0];
  _RAND_145 = {1{`RANDOM}};
  _T_1_145 = _RAND_145[20:0];
  _RAND_146 = {1{`RANDOM}};
  _T_1_146 = _RAND_146[20:0];
  _RAND_147 = {1{`RANDOM}};
  _T_1_147 = _RAND_147[20:0];
  _RAND_148 = {1{`RANDOM}};
  _T_1_148 = _RAND_148[20:0];
  _RAND_149 = {1{`RANDOM}};
  _T_1_149 = _RAND_149[20:0];
  _RAND_150 = {1{`RANDOM}};
  _T_1_150 = _RAND_150[20:0];
  _RAND_151 = {1{`RANDOM}};
  _T_1_151 = _RAND_151[20:0];
  _RAND_152 = {1{`RANDOM}};
  _T_1_152 = _RAND_152[20:0];
  _RAND_153 = {1{`RANDOM}};
  _T_1_153 = _RAND_153[20:0];
  _RAND_154 = {1{`RANDOM}};
  _T_1_154 = _RAND_154[20:0];
  _RAND_155 = {1{`RANDOM}};
  _T_1_155 = _RAND_155[20:0];
  _RAND_156 = {1{`RANDOM}};
  _T_1_156 = _RAND_156[20:0];
  _RAND_157 = {1{`RANDOM}};
  _T_1_157 = _RAND_157[20:0];
  _RAND_158 = {1{`RANDOM}};
  _T_1_158 = _RAND_158[20:0];
  _RAND_159 = {1{`RANDOM}};
  _T_1_159 = _RAND_159[20:0];
  _RAND_160 = {1{`RANDOM}};
  _T_1_160 = _RAND_160[20:0];
  _RAND_161 = {1{`RANDOM}};
  _T_1_161 = _RAND_161[20:0];
  _RAND_162 = {1{`RANDOM}};
  _T_1_162 = _RAND_162[20:0];
  _RAND_163 = {1{`RANDOM}};
  _T_1_163 = _RAND_163[20:0];
  _RAND_164 = {1{`RANDOM}};
  _T_1_164 = _RAND_164[20:0];
  _RAND_165 = {1{`RANDOM}};
  _T_1_165 = _RAND_165[20:0];
  _RAND_166 = {1{`RANDOM}};
  _T_1_166 = _RAND_166[20:0];
  _RAND_167 = {1{`RANDOM}};
  _T_1_167 = _RAND_167[20:0];
  _RAND_168 = {1{`RANDOM}};
  _T_1_168 = _RAND_168[20:0];
  _RAND_169 = {1{`RANDOM}};
  _T_1_169 = _RAND_169[20:0];
  _RAND_170 = {1{`RANDOM}};
  _T_1_170 = _RAND_170[20:0];
  _RAND_171 = {1{`RANDOM}};
  _T_1_171 = _RAND_171[20:0];
  _RAND_172 = {1{`RANDOM}};
  _T_1_172 = _RAND_172[20:0];
  _RAND_173 = {1{`RANDOM}};
  _T_1_173 = _RAND_173[20:0];
  _RAND_174 = {1{`RANDOM}};
  _T_1_174 = _RAND_174[20:0];
  _RAND_175 = {1{`RANDOM}};
  _T_1_175 = _RAND_175[20:0];
  _RAND_176 = {1{`RANDOM}};
  _T_1_176 = _RAND_176[20:0];
  _RAND_177 = {1{`RANDOM}};
  _T_1_177 = _RAND_177[20:0];
  _RAND_178 = {1{`RANDOM}};
  _T_1_178 = _RAND_178[20:0];
  _RAND_179 = {1{`RANDOM}};
  _T_1_179 = _RAND_179[20:0];
  _RAND_180 = {1{`RANDOM}};
  _T_1_180 = _RAND_180[20:0];
  _RAND_181 = {1{`RANDOM}};
  _T_1_181 = _RAND_181[20:0];
  _RAND_182 = {1{`RANDOM}};
  _T_1_182 = _RAND_182[20:0];
  _RAND_183 = {1{`RANDOM}};
  _T_1_183 = _RAND_183[20:0];
  _RAND_184 = {1{`RANDOM}};
  _T_1_184 = _RAND_184[20:0];
  _RAND_185 = {1{`RANDOM}};
  _T_1_185 = _RAND_185[20:0];
  _RAND_186 = {1{`RANDOM}};
  _T_1_186 = _RAND_186[20:0];
  _RAND_187 = {1{`RANDOM}};
  _T_1_187 = _RAND_187[20:0];
  _RAND_188 = {1{`RANDOM}};
  _T_1_188 = _RAND_188[20:0];
  _RAND_189 = {1{`RANDOM}};
  _T_1_189 = _RAND_189[20:0];
  _RAND_190 = {1{`RANDOM}};
  _T_1_190 = _RAND_190[20:0];
  _RAND_191 = {1{`RANDOM}};
  _T_1_191 = _RAND_191[20:0];
  _RAND_192 = {1{`RANDOM}};
  _T_1_192 = _RAND_192[20:0];
  _RAND_193 = {1{`RANDOM}};
  _T_1_193 = _RAND_193[20:0];
  _RAND_194 = {1{`RANDOM}};
  _T_1_194 = _RAND_194[20:0];
  _RAND_195 = {1{`RANDOM}};
  _T_1_195 = _RAND_195[20:0];
  _RAND_196 = {1{`RANDOM}};
  _T_1_196 = _RAND_196[20:0];
  _RAND_197 = {1{`RANDOM}};
  _T_1_197 = _RAND_197[20:0];
  _RAND_198 = {1{`RANDOM}};
  _T_1_198 = _RAND_198[20:0];
  _RAND_199 = {1{`RANDOM}};
  _T_1_199 = _RAND_199[20:0];
  _RAND_200 = {1{`RANDOM}};
  _T_1_200 = _RAND_200[20:0];
  _RAND_201 = {1{`RANDOM}};
  _T_1_201 = _RAND_201[20:0];
  _RAND_202 = {1{`RANDOM}};
  _T_1_202 = _RAND_202[20:0];
  _RAND_203 = {1{`RANDOM}};
  _T_1_203 = _RAND_203[20:0];
  _RAND_204 = {1{`RANDOM}};
  _T_1_204 = _RAND_204[20:0];
  _RAND_205 = {1{`RANDOM}};
  _T_1_205 = _RAND_205[20:0];
  _RAND_206 = {1{`RANDOM}};
  _T_1_206 = _RAND_206[20:0];
  _RAND_207 = {1{`RANDOM}};
  _T_1_207 = _RAND_207[20:0];
  _RAND_208 = {1{`RANDOM}};
  _T_1_208 = _RAND_208[20:0];
  _RAND_209 = {1{`RANDOM}};
  _T_1_209 = _RAND_209[20:0];
  _RAND_210 = {1{`RANDOM}};
  _T_1_210 = _RAND_210[20:0];
  _RAND_211 = {1{`RANDOM}};
  _T_1_211 = _RAND_211[20:0];
  _RAND_212 = {1{`RANDOM}};
  _T_1_212 = _RAND_212[20:0];
  _RAND_213 = {1{`RANDOM}};
  _T_1_213 = _RAND_213[20:0];
  _RAND_214 = {1{`RANDOM}};
  _T_1_214 = _RAND_214[20:0];
  _RAND_215 = {1{`RANDOM}};
  _T_1_215 = _RAND_215[20:0];
  _RAND_216 = {1{`RANDOM}};
  _T_1_216 = _RAND_216[20:0];
  _RAND_217 = {1{`RANDOM}};
  _T_1_217 = _RAND_217[20:0];
  _RAND_218 = {1{`RANDOM}};
  _T_1_218 = _RAND_218[20:0];
  _RAND_219 = {1{`RANDOM}};
  _T_1_219 = _RAND_219[20:0];
  _RAND_220 = {1{`RANDOM}};
  _T_1_220 = _RAND_220[20:0];
  _RAND_221 = {1{`RANDOM}};
  _T_1_221 = _RAND_221[20:0];
  _RAND_222 = {1{`RANDOM}};
  _T_1_222 = _RAND_222[20:0];
  _RAND_223 = {1{`RANDOM}};
  _T_1_223 = _RAND_223[20:0];
  _RAND_224 = {1{`RANDOM}};
  _T_1_224 = _RAND_224[20:0];
  _RAND_225 = {1{`RANDOM}};
  _T_1_225 = _RAND_225[20:0];
  _RAND_226 = {1{`RANDOM}};
  _T_1_226 = _RAND_226[20:0];
  _RAND_227 = {1{`RANDOM}};
  _T_1_227 = _RAND_227[20:0];
  _RAND_228 = {1{`RANDOM}};
  _T_1_228 = _RAND_228[20:0];
  _RAND_229 = {1{`RANDOM}};
  _T_1_229 = _RAND_229[20:0];
  _RAND_230 = {1{`RANDOM}};
  _T_1_230 = _RAND_230[20:0];
  _RAND_231 = {1{`RANDOM}};
  _T_1_231 = _RAND_231[20:0];
  _RAND_232 = {1{`RANDOM}};
  _T_1_232 = _RAND_232[20:0];
  _RAND_233 = {1{`RANDOM}};
  _T_1_233 = _RAND_233[20:0];
  _RAND_234 = {1{`RANDOM}};
  _T_1_234 = _RAND_234[20:0];
  _RAND_235 = {1{`RANDOM}};
  _T_1_235 = _RAND_235[20:0];
  _RAND_236 = {1{`RANDOM}};
  _T_1_236 = _RAND_236[20:0];
  _RAND_237 = {1{`RANDOM}};
  _T_1_237 = _RAND_237[20:0];
  _RAND_238 = {1{`RANDOM}};
  _T_1_238 = _RAND_238[20:0];
  _RAND_239 = {1{`RANDOM}};
  _T_1_239 = _RAND_239[20:0];
  _RAND_240 = {1{`RANDOM}};
  _T_1_240 = _RAND_240[20:0];
  _RAND_241 = {1{`RANDOM}};
  _T_1_241 = _RAND_241[20:0];
  _RAND_242 = {1{`RANDOM}};
  _T_1_242 = _RAND_242[20:0];
  _RAND_243 = {1{`RANDOM}};
  _T_1_243 = _RAND_243[20:0];
  _RAND_244 = {1{`RANDOM}};
  _T_1_244 = _RAND_244[20:0];
  _RAND_245 = {1{`RANDOM}};
  _T_1_245 = _RAND_245[20:0];
  _RAND_246 = {1{`RANDOM}};
  _T_1_246 = _RAND_246[20:0];
  _RAND_247 = {1{`RANDOM}};
  _T_1_247 = _RAND_247[20:0];
  _RAND_248 = {1{`RANDOM}};
  _T_1_248 = _RAND_248[20:0];
  _RAND_249 = {1{`RANDOM}};
  _T_1_249 = _RAND_249[20:0];
  _RAND_250 = {1{`RANDOM}};
  _T_1_250 = _RAND_250[20:0];
  _RAND_251 = {1{`RANDOM}};
  _T_1_251 = _RAND_251[20:0];
  _RAND_252 = {1{`RANDOM}};
  _T_1_252 = _RAND_252[20:0];
  _RAND_253 = {1{`RANDOM}};
  _T_1_253 = _RAND_253[20:0];
  _RAND_254 = {1{`RANDOM}};
  _T_1_254 = _RAND_254[20:0];
  _RAND_255 = {1{`RANDOM}};
  _T_1_255 = _RAND_255[20:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      _T_1_0 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h0 == io_writeAddr) begin
        _T_1_0 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_1 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h1 == io_writeAddr) begin
        _T_1_1 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_2 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h2 == io_writeAddr) begin
        _T_1_2 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_3 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h3 == io_writeAddr) begin
        _T_1_3 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_4 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h4 == io_writeAddr) begin
        _T_1_4 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_5 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h5 == io_writeAddr) begin
        _T_1_5 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_6 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h6 == io_writeAddr) begin
        _T_1_6 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_7 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h7 == io_writeAddr) begin
        _T_1_7 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_8 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h8 == io_writeAddr) begin
        _T_1_8 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_9 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h9 == io_writeAddr) begin
        _T_1_9 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_10 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'ha == io_writeAddr) begin
        _T_1_10 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_11 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'hb == io_writeAddr) begin
        _T_1_11 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_12 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'hc == io_writeAddr) begin
        _T_1_12 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_13 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'hd == io_writeAddr) begin
        _T_1_13 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_14 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'he == io_writeAddr) begin
        _T_1_14 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_15 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'hf == io_writeAddr) begin
        _T_1_15 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_16 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h10 == io_writeAddr) begin
        _T_1_16 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_17 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h11 == io_writeAddr) begin
        _T_1_17 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_18 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h12 == io_writeAddr) begin
        _T_1_18 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_19 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h13 == io_writeAddr) begin
        _T_1_19 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_20 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h14 == io_writeAddr) begin
        _T_1_20 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_21 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h15 == io_writeAddr) begin
        _T_1_21 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_22 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h16 == io_writeAddr) begin
        _T_1_22 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_23 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h17 == io_writeAddr) begin
        _T_1_23 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_24 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h18 == io_writeAddr) begin
        _T_1_24 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_25 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h19 == io_writeAddr) begin
        _T_1_25 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_26 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h1a == io_writeAddr) begin
        _T_1_26 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_27 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h1b == io_writeAddr) begin
        _T_1_27 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_28 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h1c == io_writeAddr) begin
        _T_1_28 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_29 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h1d == io_writeAddr) begin
        _T_1_29 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_30 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h1e == io_writeAddr) begin
        _T_1_30 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_31 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h1f == io_writeAddr) begin
        _T_1_31 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_32 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h20 == io_writeAddr) begin
        _T_1_32 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_33 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h21 == io_writeAddr) begin
        _T_1_33 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_34 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h22 == io_writeAddr) begin
        _T_1_34 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_35 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h23 == io_writeAddr) begin
        _T_1_35 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_36 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h24 == io_writeAddr) begin
        _T_1_36 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_37 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h25 == io_writeAddr) begin
        _T_1_37 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_38 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h26 == io_writeAddr) begin
        _T_1_38 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_39 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h27 == io_writeAddr) begin
        _T_1_39 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_40 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h28 == io_writeAddr) begin
        _T_1_40 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_41 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h29 == io_writeAddr) begin
        _T_1_41 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_42 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h2a == io_writeAddr) begin
        _T_1_42 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_43 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h2b == io_writeAddr) begin
        _T_1_43 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_44 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h2c == io_writeAddr) begin
        _T_1_44 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_45 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h2d == io_writeAddr) begin
        _T_1_45 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_46 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h2e == io_writeAddr) begin
        _T_1_46 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_47 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h2f == io_writeAddr) begin
        _T_1_47 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_48 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h30 == io_writeAddr) begin
        _T_1_48 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_49 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h31 == io_writeAddr) begin
        _T_1_49 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_50 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h32 == io_writeAddr) begin
        _T_1_50 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_51 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h33 == io_writeAddr) begin
        _T_1_51 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_52 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h34 == io_writeAddr) begin
        _T_1_52 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_53 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h35 == io_writeAddr) begin
        _T_1_53 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_54 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h36 == io_writeAddr) begin
        _T_1_54 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_55 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h37 == io_writeAddr) begin
        _T_1_55 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_56 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h38 == io_writeAddr) begin
        _T_1_56 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_57 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h39 == io_writeAddr) begin
        _T_1_57 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_58 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h3a == io_writeAddr) begin
        _T_1_58 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_59 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h3b == io_writeAddr) begin
        _T_1_59 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_60 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h3c == io_writeAddr) begin
        _T_1_60 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_61 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h3d == io_writeAddr) begin
        _T_1_61 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_62 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h3e == io_writeAddr) begin
        _T_1_62 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_63 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h3f == io_writeAddr) begin
        _T_1_63 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_64 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h40 == io_writeAddr) begin
        _T_1_64 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_65 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h41 == io_writeAddr) begin
        _T_1_65 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_66 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h42 == io_writeAddr) begin
        _T_1_66 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_67 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h43 == io_writeAddr) begin
        _T_1_67 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_68 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h44 == io_writeAddr) begin
        _T_1_68 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_69 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h45 == io_writeAddr) begin
        _T_1_69 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_70 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h46 == io_writeAddr) begin
        _T_1_70 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_71 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h47 == io_writeAddr) begin
        _T_1_71 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_72 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h48 == io_writeAddr) begin
        _T_1_72 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_73 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h49 == io_writeAddr) begin
        _T_1_73 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_74 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h4a == io_writeAddr) begin
        _T_1_74 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_75 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h4b == io_writeAddr) begin
        _T_1_75 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_76 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h4c == io_writeAddr) begin
        _T_1_76 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_77 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h4d == io_writeAddr) begin
        _T_1_77 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_78 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h4e == io_writeAddr) begin
        _T_1_78 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_79 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h4f == io_writeAddr) begin
        _T_1_79 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_80 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h50 == io_writeAddr) begin
        _T_1_80 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_81 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h51 == io_writeAddr) begin
        _T_1_81 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_82 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h52 == io_writeAddr) begin
        _T_1_82 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_83 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h53 == io_writeAddr) begin
        _T_1_83 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_84 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h54 == io_writeAddr) begin
        _T_1_84 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_85 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h55 == io_writeAddr) begin
        _T_1_85 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_86 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h56 == io_writeAddr) begin
        _T_1_86 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_87 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h57 == io_writeAddr) begin
        _T_1_87 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_88 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h58 == io_writeAddr) begin
        _T_1_88 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_89 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h59 == io_writeAddr) begin
        _T_1_89 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_90 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h5a == io_writeAddr) begin
        _T_1_90 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_91 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h5b == io_writeAddr) begin
        _T_1_91 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_92 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h5c == io_writeAddr) begin
        _T_1_92 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_93 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h5d == io_writeAddr) begin
        _T_1_93 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_94 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h5e == io_writeAddr) begin
        _T_1_94 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_95 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h5f == io_writeAddr) begin
        _T_1_95 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_96 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h60 == io_writeAddr) begin
        _T_1_96 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_97 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h61 == io_writeAddr) begin
        _T_1_97 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_98 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h62 == io_writeAddr) begin
        _T_1_98 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_99 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h63 == io_writeAddr) begin
        _T_1_99 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_100 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h64 == io_writeAddr) begin
        _T_1_100 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_101 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h65 == io_writeAddr) begin
        _T_1_101 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_102 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h66 == io_writeAddr) begin
        _T_1_102 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_103 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h67 == io_writeAddr) begin
        _T_1_103 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_104 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h68 == io_writeAddr) begin
        _T_1_104 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_105 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h69 == io_writeAddr) begin
        _T_1_105 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_106 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h6a == io_writeAddr) begin
        _T_1_106 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_107 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h6b == io_writeAddr) begin
        _T_1_107 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_108 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h6c == io_writeAddr) begin
        _T_1_108 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_109 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h6d == io_writeAddr) begin
        _T_1_109 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_110 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h6e == io_writeAddr) begin
        _T_1_110 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_111 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h6f == io_writeAddr) begin
        _T_1_111 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_112 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h70 == io_writeAddr) begin
        _T_1_112 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_113 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h71 == io_writeAddr) begin
        _T_1_113 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_114 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h72 == io_writeAddr) begin
        _T_1_114 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_115 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h73 == io_writeAddr) begin
        _T_1_115 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_116 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h74 == io_writeAddr) begin
        _T_1_116 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_117 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h75 == io_writeAddr) begin
        _T_1_117 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_118 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h76 == io_writeAddr) begin
        _T_1_118 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_119 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h77 == io_writeAddr) begin
        _T_1_119 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_120 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h78 == io_writeAddr) begin
        _T_1_120 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_121 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h79 == io_writeAddr) begin
        _T_1_121 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_122 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h7a == io_writeAddr) begin
        _T_1_122 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_123 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h7b == io_writeAddr) begin
        _T_1_123 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_124 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h7c == io_writeAddr) begin
        _T_1_124 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_125 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h7d == io_writeAddr) begin
        _T_1_125 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_126 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h7e == io_writeAddr) begin
        _T_1_126 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_127 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h7f == io_writeAddr) begin
        _T_1_127 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_128 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h80 == io_writeAddr) begin
        _T_1_128 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_129 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h81 == io_writeAddr) begin
        _T_1_129 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_130 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h82 == io_writeAddr) begin
        _T_1_130 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_131 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h83 == io_writeAddr) begin
        _T_1_131 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_132 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h84 == io_writeAddr) begin
        _T_1_132 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_133 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h85 == io_writeAddr) begin
        _T_1_133 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_134 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h86 == io_writeAddr) begin
        _T_1_134 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_135 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h87 == io_writeAddr) begin
        _T_1_135 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_136 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h88 == io_writeAddr) begin
        _T_1_136 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_137 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h89 == io_writeAddr) begin
        _T_1_137 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_138 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h8a == io_writeAddr) begin
        _T_1_138 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_139 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h8b == io_writeAddr) begin
        _T_1_139 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_140 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h8c == io_writeAddr) begin
        _T_1_140 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_141 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h8d == io_writeAddr) begin
        _T_1_141 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_142 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h8e == io_writeAddr) begin
        _T_1_142 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_143 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h8f == io_writeAddr) begin
        _T_1_143 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_144 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h90 == io_writeAddr) begin
        _T_1_144 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_145 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h91 == io_writeAddr) begin
        _T_1_145 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_146 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h92 == io_writeAddr) begin
        _T_1_146 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_147 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h93 == io_writeAddr) begin
        _T_1_147 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_148 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h94 == io_writeAddr) begin
        _T_1_148 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_149 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h95 == io_writeAddr) begin
        _T_1_149 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_150 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h96 == io_writeAddr) begin
        _T_1_150 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_151 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h97 == io_writeAddr) begin
        _T_1_151 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_152 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h98 == io_writeAddr) begin
        _T_1_152 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_153 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h99 == io_writeAddr) begin
        _T_1_153 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_154 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h9a == io_writeAddr) begin
        _T_1_154 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_155 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h9b == io_writeAddr) begin
        _T_1_155 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_156 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h9c == io_writeAddr) begin
        _T_1_156 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_157 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h9d == io_writeAddr) begin
        _T_1_157 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_158 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h9e == io_writeAddr) begin
        _T_1_158 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_159 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'h9f == io_writeAddr) begin
        _T_1_159 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_160 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'ha0 == io_writeAddr) begin
        _T_1_160 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_161 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'ha1 == io_writeAddr) begin
        _T_1_161 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_162 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'ha2 == io_writeAddr) begin
        _T_1_162 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_163 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'ha3 == io_writeAddr) begin
        _T_1_163 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_164 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'ha4 == io_writeAddr) begin
        _T_1_164 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_165 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'ha5 == io_writeAddr) begin
        _T_1_165 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_166 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'ha6 == io_writeAddr) begin
        _T_1_166 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_167 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'ha7 == io_writeAddr) begin
        _T_1_167 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_168 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'ha8 == io_writeAddr) begin
        _T_1_168 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_169 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'ha9 == io_writeAddr) begin
        _T_1_169 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_170 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'haa == io_writeAddr) begin
        _T_1_170 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_171 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'hab == io_writeAddr) begin
        _T_1_171 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_172 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'hac == io_writeAddr) begin
        _T_1_172 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_173 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'had == io_writeAddr) begin
        _T_1_173 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_174 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'hae == io_writeAddr) begin
        _T_1_174 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_175 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'haf == io_writeAddr) begin
        _T_1_175 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_176 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'hb0 == io_writeAddr) begin
        _T_1_176 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_177 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'hb1 == io_writeAddr) begin
        _T_1_177 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_178 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'hb2 == io_writeAddr) begin
        _T_1_178 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_179 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'hb3 == io_writeAddr) begin
        _T_1_179 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_180 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'hb4 == io_writeAddr) begin
        _T_1_180 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_181 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'hb5 == io_writeAddr) begin
        _T_1_181 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_182 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'hb6 == io_writeAddr) begin
        _T_1_182 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_183 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'hb7 == io_writeAddr) begin
        _T_1_183 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_184 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'hb8 == io_writeAddr) begin
        _T_1_184 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_185 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'hb9 == io_writeAddr) begin
        _T_1_185 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_186 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'hba == io_writeAddr) begin
        _T_1_186 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_187 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'hbb == io_writeAddr) begin
        _T_1_187 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_188 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'hbc == io_writeAddr) begin
        _T_1_188 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_189 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'hbd == io_writeAddr) begin
        _T_1_189 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_190 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'hbe == io_writeAddr) begin
        _T_1_190 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_191 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'hbf == io_writeAddr) begin
        _T_1_191 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_192 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'hc0 == io_writeAddr) begin
        _T_1_192 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_193 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'hc1 == io_writeAddr) begin
        _T_1_193 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_194 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'hc2 == io_writeAddr) begin
        _T_1_194 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_195 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'hc3 == io_writeAddr) begin
        _T_1_195 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_196 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'hc4 == io_writeAddr) begin
        _T_1_196 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_197 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'hc5 == io_writeAddr) begin
        _T_1_197 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_198 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'hc6 == io_writeAddr) begin
        _T_1_198 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_199 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'hc7 == io_writeAddr) begin
        _T_1_199 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_200 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'hc8 == io_writeAddr) begin
        _T_1_200 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_201 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'hc9 == io_writeAddr) begin
        _T_1_201 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_202 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'hca == io_writeAddr) begin
        _T_1_202 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_203 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'hcb == io_writeAddr) begin
        _T_1_203 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_204 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'hcc == io_writeAddr) begin
        _T_1_204 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_205 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'hcd == io_writeAddr) begin
        _T_1_205 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_206 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'hce == io_writeAddr) begin
        _T_1_206 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_207 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'hcf == io_writeAddr) begin
        _T_1_207 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_208 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'hd0 == io_writeAddr) begin
        _T_1_208 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_209 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'hd1 == io_writeAddr) begin
        _T_1_209 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_210 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'hd2 == io_writeAddr) begin
        _T_1_210 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_211 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'hd3 == io_writeAddr) begin
        _T_1_211 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_212 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'hd4 == io_writeAddr) begin
        _T_1_212 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_213 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'hd5 == io_writeAddr) begin
        _T_1_213 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_214 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'hd6 == io_writeAddr) begin
        _T_1_214 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_215 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'hd7 == io_writeAddr) begin
        _T_1_215 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_216 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'hd8 == io_writeAddr) begin
        _T_1_216 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_217 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'hd9 == io_writeAddr) begin
        _T_1_217 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_218 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'hda == io_writeAddr) begin
        _T_1_218 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_219 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'hdb == io_writeAddr) begin
        _T_1_219 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_220 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'hdc == io_writeAddr) begin
        _T_1_220 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_221 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'hdd == io_writeAddr) begin
        _T_1_221 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_222 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'hde == io_writeAddr) begin
        _T_1_222 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_223 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'hdf == io_writeAddr) begin
        _T_1_223 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_224 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'he0 == io_writeAddr) begin
        _T_1_224 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_225 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'he1 == io_writeAddr) begin
        _T_1_225 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_226 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'he2 == io_writeAddr) begin
        _T_1_226 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_227 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'he3 == io_writeAddr) begin
        _T_1_227 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_228 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'he4 == io_writeAddr) begin
        _T_1_228 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_229 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'he5 == io_writeAddr) begin
        _T_1_229 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_230 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'he6 == io_writeAddr) begin
        _T_1_230 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_231 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'he7 == io_writeAddr) begin
        _T_1_231 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_232 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'he8 == io_writeAddr) begin
        _T_1_232 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_233 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'he9 == io_writeAddr) begin
        _T_1_233 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_234 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'hea == io_writeAddr) begin
        _T_1_234 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_235 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'heb == io_writeAddr) begin
        _T_1_235 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_236 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'hec == io_writeAddr) begin
        _T_1_236 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_237 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'hed == io_writeAddr) begin
        _T_1_237 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_238 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'hee == io_writeAddr) begin
        _T_1_238 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_239 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'hef == io_writeAddr) begin
        _T_1_239 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_240 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'hf0 == io_writeAddr) begin
        _T_1_240 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_241 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'hf1 == io_writeAddr) begin
        _T_1_241 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_242 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'hf2 == io_writeAddr) begin
        _T_1_242 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_243 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'hf3 == io_writeAddr) begin
        _T_1_243 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_244 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'hf4 == io_writeAddr) begin
        _T_1_244 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_245 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'hf5 == io_writeAddr) begin
        _T_1_245 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_246 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'hf6 == io_writeAddr) begin
        _T_1_246 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_247 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'hf7 == io_writeAddr) begin
        _T_1_247 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_248 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'hf8 == io_writeAddr) begin
        _T_1_248 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_249 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'hf9 == io_writeAddr) begin
        _T_1_249 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_250 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'hfa == io_writeAddr) begin
        _T_1_250 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_251 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'hfb == io_writeAddr) begin
        _T_1_251 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_252 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'hfc == io_writeAddr) begin
        _T_1_252 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_253 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'hfd == io_writeAddr) begin
        _T_1_253 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_254 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'hfe == io_writeAddr) begin
        _T_1_254 <= io_writeData;
      end
    end
    if (reset) begin
      _T_1_255 <= 21'h0;
    end else if (io_writeEnable) begin
      if (8'hff == io_writeAddr) begin
        _T_1_255 <= io_writeData;
      end
    end
  end
endmodule
module TagValidBanks(
  input         clock,
  input         reset,
  input  [7:0]  io_way_0_portA_addr,
  output [19:0] io_way_0_portA_data_tag,
  output        io_way_0_portA_data_valid,
  input  [7:0]  io_way_0_portB_addr,
  input         io_way_0_portB_writeEnable,
  input  [19:0] io_way_0_portB_writeData_tag,
  input  [7:0]  io_way_1_portA_addr,
  output [19:0] io_way_1_portA_data_tag,
  output        io_way_1_portA_data_valid,
  input  [7:0]  io_way_1_portB_addr,
  input         io_way_1_portB_writeEnable,
  input  [19:0] io_way_1_portB_writeData_tag,
  input  [7:0]  io_way_2_portA_addr,
  output [19:0] io_way_2_portA_data_tag,
  output        io_way_2_portA_data_valid,
  input  [7:0]  io_way_2_portB_addr,
  input         io_way_2_portB_writeEnable,
  input  [19:0] io_way_2_portB_writeData_tag,
  input  [7:0]  io_way_3_portA_addr,
  output [19:0] io_way_3_portA_data_tag,
  output        io_way_3_portA_data_valid,
  input  [7:0]  io_way_3_portB_addr,
  input         io_way_3_portB_writeEnable,
  input  [19:0] io_way_3_portB_writeData_tag
);
  wire  tag_valid_bank_way_0_clock; // @[TagValidBanks.scala 53:22]
  wire  tag_valid_bank_way_0_reset; // @[TagValidBanks.scala 53:22]
  wire [7:0] tag_valid_bank_way_0_io_readAddr; // @[TagValidBanks.scala 53:22]
  wire [20:0] tag_valid_bank_way_0_io_readData; // @[TagValidBanks.scala 53:22]
  wire [7:0] tag_valid_bank_way_0_io_writeAddr; // @[TagValidBanks.scala 53:22]
  wire [20:0] tag_valid_bank_way_0_io_writeData; // @[TagValidBanks.scala 53:22]
  wire  tag_valid_bank_way_0_io_writeEnable; // @[TagValidBanks.scala 53:22]
  wire  tag_valid_bank_way_1_clock; // @[TagValidBanks.scala 53:22]
  wire  tag_valid_bank_way_1_reset; // @[TagValidBanks.scala 53:22]
  wire [7:0] tag_valid_bank_way_1_io_readAddr; // @[TagValidBanks.scala 53:22]
  wire [20:0] tag_valid_bank_way_1_io_readData; // @[TagValidBanks.scala 53:22]
  wire [7:0] tag_valid_bank_way_1_io_writeAddr; // @[TagValidBanks.scala 53:22]
  wire [20:0] tag_valid_bank_way_1_io_writeData; // @[TagValidBanks.scala 53:22]
  wire  tag_valid_bank_way_1_io_writeEnable; // @[TagValidBanks.scala 53:22]
  wire  tag_valid_bank_way_2_clock; // @[TagValidBanks.scala 53:22]
  wire  tag_valid_bank_way_2_reset; // @[TagValidBanks.scala 53:22]
  wire [7:0] tag_valid_bank_way_2_io_readAddr; // @[TagValidBanks.scala 53:22]
  wire [20:0] tag_valid_bank_way_2_io_readData; // @[TagValidBanks.scala 53:22]
  wire [7:0] tag_valid_bank_way_2_io_writeAddr; // @[TagValidBanks.scala 53:22]
  wire [20:0] tag_valid_bank_way_2_io_writeData; // @[TagValidBanks.scala 53:22]
  wire  tag_valid_bank_way_2_io_writeEnable; // @[TagValidBanks.scala 53:22]
  wire  tag_valid_bank_way_3_clock; // @[TagValidBanks.scala 53:22]
  wire  tag_valid_bank_way_3_reset; // @[TagValidBanks.scala 53:22]
  wire [7:0] tag_valid_bank_way_3_io_readAddr; // @[TagValidBanks.scala 53:22]
  wire [20:0] tag_valid_bank_way_3_io_readData; // @[TagValidBanks.scala 53:22]
  wire [7:0] tag_valid_bank_way_3_io_writeAddr; // @[TagValidBanks.scala 53:22]
  wire [20:0] tag_valid_bank_way_3_io_writeData; // @[TagValidBanks.scala 53:22]
  wire  tag_valid_bank_way_3_io_writeEnable; // @[TagValidBanks.scala 53:22]
  wire [20:0] _T_1 = tag_valid_bank_way_0_io_readData;
  wire [20:0] _T_11 = tag_valid_bank_way_1_io_readData;
  wire [20:0] _T_21 = tag_valid_bank_way_2_io_readData;
  wire [20:0] _T_31 = tag_valid_bank_way_3_io_readData;
  LUTRam tag_valid_bank_way_0 ( // @[TagValidBanks.scala 53:22]
    .clock(tag_valid_bank_way_0_clock),
    .reset(tag_valid_bank_way_0_reset),
    .io_readAddr(tag_valid_bank_way_0_io_readAddr),
    .io_readData(tag_valid_bank_way_0_io_readData),
    .io_writeAddr(tag_valid_bank_way_0_io_writeAddr),
    .io_writeData(tag_valid_bank_way_0_io_writeData),
    .io_writeEnable(tag_valid_bank_way_0_io_writeEnable)
  );
  LUTRam tag_valid_bank_way_1 ( // @[TagValidBanks.scala 53:22]
    .clock(tag_valid_bank_way_1_clock),
    .reset(tag_valid_bank_way_1_reset),
    .io_readAddr(tag_valid_bank_way_1_io_readAddr),
    .io_readData(tag_valid_bank_way_1_io_readData),
    .io_writeAddr(tag_valid_bank_way_1_io_writeAddr),
    .io_writeData(tag_valid_bank_way_1_io_writeData),
    .io_writeEnable(tag_valid_bank_way_1_io_writeEnable)
  );
  LUTRam tag_valid_bank_way_2 ( // @[TagValidBanks.scala 53:22]
    .clock(tag_valid_bank_way_2_clock),
    .reset(tag_valid_bank_way_2_reset),
    .io_readAddr(tag_valid_bank_way_2_io_readAddr),
    .io_readData(tag_valid_bank_way_2_io_readData),
    .io_writeAddr(tag_valid_bank_way_2_io_writeAddr),
    .io_writeData(tag_valid_bank_way_2_io_writeData),
    .io_writeEnable(tag_valid_bank_way_2_io_writeEnable)
  );
  LUTRam tag_valid_bank_way_3 ( // @[TagValidBanks.scala 53:22]
    .clock(tag_valid_bank_way_3_clock),
    .reset(tag_valid_bank_way_3_reset),
    .io_readAddr(tag_valid_bank_way_3_io_readAddr),
    .io_readData(tag_valid_bank_way_3_io_readData),
    .io_writeAddr(tag_valid_bank_way_3_io_writeAddr),
    .io_writeData(tag_valid_bank_way_3_io_writeData),
    .io_writeEnable(tag_valid_bank_way_3_io_writeEnable)
  );
  assign io_way_0_portA_data_tag = _T_1[20:1]; // @[TagValidBanks.scala 56:26]
  assign io_way_0_portA_data_valid = _T_1[0]; // @[TagValidBanks.scala 56:26]
  assign io_way_1_portA_data_tag = _T_11[20:1]; // @[TagValidBanks.scala 56:26]
  assign io_way_1_portA_data_valid = _T_11[0]; // @[TagValidBanks.scala 56:26]
  assign io_way_2_portA_data_tag = _T_21[20:1]; // @[TagValidBanks.scala 56:26]
  assign io_way_2_portA_data_valid = _T_21[0]; // @[TagValidBanks.scala 56:26]
  assign io_way_3_portA_data_tag = _T_31[20:1]; // @[TagValidBanks.scala 56:26]
  assign io_way_3_portA_data_valid = _T_31[0]; // @[TagValidBanks.scala 56:26]
  assign tag_valid_bank_way_0_clock = clock;
  assign tag_valid_bank_way_0_reset = reset;
  assign tag_valid_bank_way_0_io_readAddr = io_way_0_portA_addr; // @[TagValidBanks.scala 55:22]
  assign tag_valid_bank_way_0_io_writeAddr = io_way_0_portB_addr; // @[TagValidBanks.scala 58:23]
  assign tag_valid_bank_way_0_io_writeData = {io_way_0_portB_writeData_tag,1'h1}; // @[TagValidBanks.scala 60:23]
  assign tag_valid_bank_way_0_io_writeEnable = io_way_0_portB_writeEnable; // @[TagValidBanks.scala 59:25]
  assign tag_valid_bank_way_1_clock = clock;
  assign tag_valid_bank_way_1_reset = reset;
  assign tag_valid_bank_way_1_io_readAddr = io_way_1_portA_addr; // @[TagValidBanks.scala 55:22]
  assign tag_valid_bank_way_1_io_writeAddr = io_way_1_portB_addr; // @[TagValidBanks.scala 58:23]
  assign tag_valid_bank_way_1_io_writeData = {io_way_1_portB_writeData_tag,1'h1}; // @[TagValidBanks.scala 60:23]
  assign tag_valid_bank_way_1_io_writeEnable = io_way_1_portB_writeEnable; // @[TagValidBanks.scala 59:25]
  assign tag_valid_bank_way_2_clock = clock;
  assign tag_valid_bank_way_2_reset = reset;
  assign tag_valid_bank_way_2_io_readAddr = io_way_2_portA_addr; // @[TagValidBanks.scala 55:22]
  assign tag_valid_bank_way_2_io_writeAddr = io_way_2_portB_addr; // @[TagValidBanks.scala 58:23]
  assign tag_valid_bank_way_2_io_writeData = {io_way_2_portB_writeData_tag,1'h1}; // @[TagValidBanks.scala 60:23]
  assign tag_valid_bank_way_2_io_writeEnable = io_way_2_portB_writeEnable; // @[TagValidBanks.scala 59:25]
  assign tag_valid_bank_way_3_clock = clock;
  assign tag_valid_bank_way_3_reset = reset;
  assign tag_valid_bank_way_3_io_readAddr = io_way_3_portA_addr; // @[TagValidBanks.scala 55:22]
  assign tag_valid_bank_way_3_io_writeAddr = io_way_3_portB_addr; // @[TagValidBanks.scala 58:23]
  assign tag_valid_bank_way_3_io_writeData = {io_way_3_portB_writeData_tag,1'h1}; // @[TagValidBanks.scala 60:23]
  assign tag_valid_bank_way_3_io_writeEnable = io_way_3_portB_writeEnable; // @[TagValidBanks.scala 59:25]
endmodule
module TagValid(
  input         clock,
  input         reset,
  input  [7:0]  io_address,
  input         io_write_valid,
  input  [1:0]  io_write_bits_waySelection,
  input  [7:0]  io_write_bits_indexSelection,
  input  [19:0] io_write_bits_tagValid_tag,
  output [19:0] io_tagValid_0_tag,
  output        io_tagValid_0_valid,
  output [19:0] io_tagValid_1_tag,
  output        io_tagValid_1_valid,
  output [19:0] io_tagValid_2_tag,
  output        io_tagValid_2_valid,
  output [19:0] io_tagValid_3_tag,
  output        io_tagValid_3_valid
);
  wire  tagValidBanks_clock; // @[TagValid.scala 28:29]
  wire  tagValidBanks_reset; // @[TagValid.scala 28:29]
  wire [7:0] tagValidBanks_io_way_0_portA_addr; // @[TagValid.scala 28:29]
  wire [19:0] tagValidBanks_io_way_0_portA_data_tag; // @[TagValid.scala 28:29]
  wire  tagValidBanks_io_way_0_portA_data_valid; // @[TagValid.scala 28:29]
  wire [7:0] tagValidBanks_io_way_0_portB_addr; // @[TagValid.scala 28:29]
  wire  tagValidBanks_io_way_0_portB_writeEnable; // @[TagValid.scala 28:29]
  wire [19:0] tagValidBanks_io_way_0_portB_writeData_tag; // @[TagValid.scala 28:29]
  wire [7:0] tagValidBanks_io_way_1_portA_addr; // @[TagValid.scala 28:29]
  wire [19:0] tagValidBanks_io_way_1_portA_data_tag; // @[TagValid.scala 28:29]
  wire  tagValidBanks_io_way_1_portA_data_valid; // @[TagValid.scala 28:29]
  wire [7:0] tagValidBanks_io_way_1_portB_addr; // @[TagValid.scala 28:29]
  wire  tagValidBanks_io_way_1_portB_writeEnable; // @[TagValid.scala 28:29]
  wire [19:0] tagValidBanks_io_way_1_portB_writeData_tag; // @[TagValid.scala 28:29]
  wire [7:0] tagValidBanks_io_way_2_portA_addr; // @[TagValid.scala 28:29]
  wire [19:0] tagValidBanks_io_way_2_portA_data_tag; // @[TagValid.scala 28:29]
  wire  tagValidBanks_io_way_2_portA_data_valid; // @[TagValid.scala 28:29]
  wire [7:0] tagValidBanks_io_way_2_portB_addr; // @[TagValid.scala 28:29]
  wire  tagValidBanks_io_way_2_portB_writeEnable; // @[TagValid.scala 28:29]
  wire [19:0] tagValidBanks_io_way_2_portB_writeData_tag; // @[TagValid.scala 28:29]
  wire [7:0] tagValidBanks_io_way_3_portA_addr; // @[TagValid.scala 28:29]
  wire [19:0] tagValidBanks_io_way_3_portA_data_tag; // @[TagValid.scala 28:29]
  wire  tagValidBanks_io_way_3_portA_data_valid; // @[TagValid.scala 28:29]
  wire [7:0] tagValidBanks_io_way_3_portB_addr; // @[TagValid.scala 28:29]
  wire  tagValidBanks_io_way_3_portB_writeEnable; // @[TagValid.scala 28:29]
  wire [19:0] tagValidBanks_io_way_3_portB_writeData_tag; // @[TagValid.scala 28:29]
  wire  _T = io_write_bits_waySelection == 2'h0; // @[TagValid.scala 38:98]
  wire  _T_3 = io_write_bits_waySelection == 2'h1; // @[TagValid.scala 38:98]
  wire  _T_6 = io_write_bits_waySelection == 2'h2; // @[TagValid.scala 38:98]
  wire  _T_9 = io_write_bits_waySelection == 2'h3; // @[TagValid.scala 38:98]
  TagValidBanks tagValidBanks ( // @[TagValid.scala 28:29]
    .clock(tagValidBanks_clock),
    .reset(tagValidBanks_reset),
    .io_way_0_portA_addr(tagValidBanks_io_way_0_portA_addr),
    .io_way_0_portA_data_tag(tagValidBanks_io_way_0_portA_data_tag),
    .io_way_0_portA_data_valid(tagValidBanks_io_way_0_portA_data_valid),
    .io_way_0_portB_addr(tagValidBanks_io_way_0_portB_addr),
    .io_way_0_portB_writeEnable(tagValidBanks_io_way_0_portB_writeEnable),
    .io_way_0_portB_writeData_tag(tagValidBanks_io_way_0_portB_writeData_tag),
    .io_way_1_portA_addr(tagValidBanks_io_way_1_portA_addr),
    .io_way_1_portA_data_tag(tagValidBanks_io_way_1_portA_data_tag),
    .io_way_1_portA_data_valid(tagValidBanks_io_way_1_portA_data_valid),
    .io_way_1_portB_addr(tagValidBanks_io_way_1_portB_addr),
    .io_way_1_portB_writeEnable(tagValidBanks_io_way_1_portB_writeEnable),
    .io_way_1_portB_writeData_tag(tagValidBanks_io_way_1_portB_writeData_tag),
    .io_way_2_portA_addr(tagValidBanks_io_way_2_portA_addr),
    .io_way_2_portA_data_tag(tagValidBanks_io_way_2_portA_data_tag),
    .io_way_2_portA_data_valid(tagValidBanks_io_way_2_portA_data_valid),
    .io_way_2_portB_addr(tagValidBanks_io_way_2_portB_addr),
    .io_way_2_portB_writeEnable(tagValidBanks_io_way_2_portB_writeEnable),
    .io_way_2_portB_writeData_tag(tagValidBanks_io_way_2_portB_writeData_tag),
    .io_way_3_portA_addr(tagValidBanks_io_way_3_portA_addr),
    .io_way_3_portA_data_tag(tagValidBanks_io_way_3_portA_data_tag),
    .io_way_3_portA_data_valid(tagValidBanks_io_way_3_portA_data_valid),
    .io_way_3_portB_addr(tagValidBanks_io_way_3_portB_addr),
    .io_way_3_portB_writeEnable(tagValidBanks_io_way_3_portB_writeEnable),
    .io_way_3_portB_writeData_tag(tagValidBanks_io_way_3_portB_writeData_tag)
  );
  assign io_tagValid_0_tag = tagValidBanks_io_way_0_portA_data_tag; // @[TagValid.scala 34:40]
  assign io_tagValid_0_valid = tagValidBanks_io_way_0_portA_data_valid; // @[TagValid.scala 34:40]
  assign io_tagValid_1_tag = tagValidBanks_io_way_1_portA_data_tag; // @[TagValid.scala 34:40]
  assign io_tagValid_1_valid = tagValidBanks_io_way_1_portA_data_valid; // @[TagValid.scala 34:40]
  assign io_tagValid_2_tag = tagValidBanks_io_way_2_portA_data_tag; // @[TagValid.scala 34:40]
  assign io_tagValid_2_valid = tagValidBanks_io_way_2_portA_data_valid; // @[TagValid.scala 34:40]
  assign io_tagValid_3_tag = tagValidBanks_io_way_3_portA_data_tag; // @[TagValid.scala 34:40]
  assign io_tagValid_3_valid = tagValidBanks_io_way_3_portA_data_valid; // @[TagValid.scala 34:40]
  assign tagValidBanks_clock = clock;
  assign tagValidBanks_reset = reset;
  assign tagValidBanks_io_way_0_portA_addr = io_address; // @[TagValid.scala 33:40]
  assign tagValidBanks_io_way_0_portB_addr = io_write_bits_indexSelection; // @[TagValid.scala 37:49]
  assign tagValidBanks_io_way_0_portB_writeEnable = io_write_valid & _T; // @[TagValid.scala 38:49]
  assign tagValidBanks_io_way_0_portB_writeData_tag = io_write_bits_tagValid_tag; // @[TagValid.scala 39:49]
  assign tagValidBanks_io_way_1_portA_addr = io_address; // @[TagValid.scala 33:40]
  assign tagValidBanks_io_way_1_portB_addr = io_write_bits_indexSelection; // @[TagValid.scala 37:49]
  assign tagValidBanks_io_way_1_portB_writeEnable = io_write_valid & _T_3; // @[TagValid.scala 38:49]
  assign tagValidBanks_io_way_1_portB_writeData_tag = io_write_bits_tagValid_tag; // @[TagValid.scala 39:49]
  assign tagValidBanks_io_way_2_portA_addr = io_address; // @[TagValid.scala 33:40]
  assign tagValidBanks_io_way_2_portB_addr = io_write_bits_indexSelection; // @[TagValid.scala 37:49]
  assign tagValidBanks_io_way_2_portB_writeEnable = io_write_valid & _T_6; // @[TagValid.scala 38:49]
  assign tagValidBanks_io_way_2_portB_writeData_tag = io_write_bits_tagValid_tag; // @[TagValid.scala 39:49]
  assign tagValidBanks_io_way_3_portA_addr = io_address; // @[TagValid.scala 33:40]
  assign tagValidBanks_io_way_3_portB_addr = io_write_bits_indexSelection; // @[TagValid.scala 37:49]
  assign tagValidBanks_io_way_3_portB_writeEnable = io_write_valid & _T_9; // @[TagValid.scala 38:49]
  assign tagValidBanks_io_way_3_portB_writeData_tag = io_write_bits_tagValid_tag; // @[TagValid.scala 39:49]
endmodule
module FetchTop(
  input         clock,
  input         reset,
  input  [31:0] io_addr,
  input         io_writeTagValid_valid,
  input  [1:0]  io_writeTagValid_bits_waySelection,
  input  [7:0]  io_writeTagValid_bits_indexSelection,
  input  [19:0] io_writeTagValid_bits_tagValid_tag,
  output [7:0]  io_index,
  output [19:0] io_tagValid_0_tag,
  output        io_tagValid_0_valid,
  output [19:0] io_tagValid_1_tag,
  output        io_tagValid_1_valid,
  output [19:0] io_tagValid_2_tag,
  output        io_tagValid_2_valid,
  output [19:0] io_tagValid_3_tag,
  output        io_tagValid_3_valid,
  output [19:0] io_phyTag,
  output        io_bankIndex
);
  wire  tagValid_clock; // @[FetchTop.scala 32:24]
  wire  tagValid_reset; // @[FetchTop.scala 32:24]
  wire [7:0] tagValid_io_address; // @[FetchTop.scala 32:24]
  wire  tagValid_io_write_valid; // @[FetchTop.scala 32:24]
  wire [1:0] tagValid_io_write_bits_waySelection; // @[FetchTop.scala 32:24]
  wire [7:0] tagValid_io_write_bits_indexSelection; // @[FetchTop.scala 32:24]
  wire [19:0] tagValid_io_write_bits_tagValid_tag; // @[FetchTop.scala 32:24]
  wire [19:0] tagValid_io_tagValid_0_tag; // @[FetchTop.scala 32:24]
  wire  tagValid_io_tagValid_0_valid; // @[FetchTop.scala 32:24]
  wire [19:0] tagValid_io_tagValid_1_tag; // @[FetchTop.scala 32:24]
  wire  tagValid_io_tagValid_1_valid; // @[FetchTop.scala 32:24]
  wire [19:0] tagValid_io_tagValid_2_tag; // @[FetchTop.scala 32:24]
  wire  tagValid_io_tagValid_2_valid; // @[FetchTop.scala 32:24]
  wire [19:0] tagValid_io_tagValid_3_tag; // @[FetchTop.scala 32:24]
  wire  tagValid_io_tagValid_3_valid; // @[FetchTop.scala 32:24]
  wire [19:0] virtualTag = io_addr[31:12]; // @[FetchTop.scala 34:27]
  TagValid tagValid ( // @[FetchTop.scala 32:24]
    .clock(tagValid_clock),
    .reset(tagValid_reset),
    .io_address(tagValid_io_address),
    .io_write_valid(tagValid_io_write_valid),
    .io_write_bits_waySelection(tagValid_io_write_bits_waySelection),
    .io_write_bits_indexSelection(tagValid_io_write_bits_indexSelection),
    .io_write_bits_tagValid_tag(tagValid_io_write_bits_tagValid_tag),
    .io_tagValid_0_tag(tagValid_io_tagValid_0_tag),
    .io_tagValid_0_valid(tagValid_io_tagValid_0_valid),
    .io_tagValid_1_tag(tagValid_io_tagValid_1_tag),
    .io_tagValid_1_valid(tagValid_io_tagValid_1_valid),
    .io_tagValid_2_tag(tagValid_io_tagValid_2_tag),
    .io_tagValid_2_valid(tagValid_io_tagValid_2_valid),
    .io_tagValid_3_tag(tagValid_io_tagValid_3_tag),
    .io_tagValid_3_valid(tagValid_io_tagValid_3_valid)
  );
  assign io_index = io_addr[10:3]; // @[FetchTop.scala 41:23]
  assign io_tagValid_0_tag = tagValid_io_tagValid_0_tag; // @[FetchTop.scala 44:23]
  assign io_tagValid_0_valid = tagValid_io_tagValid_0_valid; // @[FetchTop.scala 44:23]
  assign io_tagValid_1_tag = tagValid_io_tagValid_1_tag; // @[FetchTop.scala 44:23]
  assign io_tagValid_1_valid = tagValid_io_tagValid_1_valid; // @[FetchTop.scala 44:23]
  assign io_tagValid_2_tag = tagValid_io_tagValid_2_tag; // @[FetchTop.scala 44:23]
  assign io_tagValid_2_valid = tagValid_io_tagValid_2_valid; // @[FetchTop.scala 44:23]
  assign io_tagValid_3_tag = tagValid_io_tagValid_3_tag; // @[FetchTop.scala 44:23]
  assign io_tagValid_3_valid = tagValid_io_tagValid_3_valid; // @[FetchTop.scala 44:23]
  assign io_phyTag = {3'h0,virtualTag[16:0]}; // @[FetchTop.scala 47:13]
  assign io_bankIndex = io_addr[2]; // @[FetchTop.scala 45:23]
  assign tagValid_clock = clock;
  assign tagValid_reset = reset;
  assign tagValid_io_address = io_addr[10:3]; // @[FetchTop.scala 42:23]
  assign tagValid_io_write_valid = io_writeTagValid_valid; // @[FetchTop.scala 43:23]
  assign tagValid_io_write_bits_waySelection = io_writeTagValid_bits_waySelection; // @[FetchTop.scala 43:23]
  assign tagValid_io_write_bits_indexSelection = io_writeTagValid_bits_indexSelection; // @[FetchTop.scala 43:23]
  assign tagValid_io_write_bits_tagValid_tag = io_writeTagValid_bits_tagValid_tag; // @[FetchTop.scala 43:23]
endmodule
module CachePipelineStage(
  input         clock,
  input         reset,
  input         io_stall,
  input  [19:0] io_in_tagValid_0_tag,
  input         io_in_tagValid_0_valid,
  input  [19:0] io_in_tagValid_1_tag,
  input         io_in_tagValid_1_valid,
  input  [19:0] io_in_tagValid_2_tag,
  input         io_in_tagValid_2_valid,
  input  [19:0] io_in_tagValid_3_tag,
  input         io_in_tagValid_3_valid,
  input  [19:0] io_in_phyTag,
  input  [7:0]  io_in_index,
  input         io_in_bankIndex,
  input         io_in_valid,
  output [19:0] io_out_tagValid_0_tag,
  output        io_out_tagValid_0_valid,
  output [19:0] io_out_tagValid_1_tag,
  output        io_out_tagValid_1_valid,
  output [19:0] io_out_tagValid_2_tag,
  output        io_out_tagValid_2_valid,
  output [19:0] io_out_tagValid_3_tag,
  output        io_out_tagValid_3_valid,
  output [19:0] io_out_phyTag,
  output [7:0]  io_out_index,
  output        io_out_bankIndex,
  output        io_out_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
`endif // RANDOMIZE_REG_INIT
  reg [19:0] pipelineReg_tagValid_0_tag; // @[CachePipelineStage.scala 24:28]
  reg  pipelineReg_tagValid_0_valid; // @[CachePipelineStage.scala 24:28]
  reg [19:0] pipelineReg_tagValid_1_tag; // @[CachePipelineStage.scala 24:28]
  reg  pipelineReg_tagValid_1_valid; // @[CachePipelineStage.scala 24:28]
  reg [19:0] pipelineReg_tagValid_2_tag; // @[CachePipelineStage.scala 24:28]
  reg  pipelineReg_tagValid_2_valid; // @[CachePipelineStage.scala 24:28]
  reg [19:0] pipelineReg_tagValid_3_tag; // @[CachePipelineStage.scala 24:28]
  reg  pipelineReg_tagValid_3_valid; // @[CachePipelineStage.scala 24:28]
  reg [19:0] pipelineReg_phyTag; // @[CachePipelineStage.scala 24:28]
  reg [7:0] pipelineReg_index; // @[CachePipelineStage.scala 24:28]
  reg  pipelineReg_bankIndex; // @[CachePipelineStage.scala 24:28]
  reg  pipelineReg_valid; // @[CachePipelineStage.scala 24:28]
  wire  _T_1 = ~io_stall; // @[CachePipelineStage.scala 26:8]
  assign io_out_tagValid_0_tag = pipelineReg_tagValid_0_tag; // @[CachePipelineStage.scala 30:10]
  assign io_out_tagValid_0_valid = pipelineReg_tagValid_0_valid; // @[CachePipelineStage.scala 30:10]
  assign io_out_tagValid_1_tag = pipelineReg_tagValid_1_tag; // @[CachePipelineStage.scala 30:10]
  assign io_out_tagValid_1_valid = pipelineReg_tagValid_1_valid; // @[CachePipelineStage.scala 30:10]
  assign io_out_tagValid_2_tag = pipelineReg_tagValid_2_tag; // @[CachePipelineStage.scala 30:10]
  assign io_out_tagValid_2_valid = pipelineReg_tagValid_2_valid; // @[CachePipelineStage.scala 30:10]
  assign io_out_tagValid_3_tag = pipelineReg_tagValid_3_tag; // @[CachePipelineStage.scala 30:10]
  assign io_out_tagValid_3_valid = pipelineReg_tagValid_3_valid; // @[CachePipelineStage.scala 30:10]
  assign io_out_phyTag = pipelineReg_phyTag; // @[CachePipelineStage.scala 30:10]
  assign io_out_index = pipelineReg_index; // @[CachePipelineStage.scala 30:10]
  assign io_out_bankIndex = pipelineReg_bankIndex; // @[CachePipelineStage.scala 30:10]
  assign io_out_valid = pipelineReg_valid; // @[CachePipelineStage.scala 30:10]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  pipelineReg_tagValid_0_tag = _RAND_0[19:0];
  _RAND_1 = {1{`RANDOM}};
  pipelineReg_tagValid_0_valid = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  pipelineReg_tagValid_1_tag = _RAND_2[19:0];
  _RAND_3 = {1{`RANDOM}};
  pipelineReg_tagValid_1_valid = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  pipelineReg_tagValid_2_tag = _RAND_4[19:0];
  _RAND_5 = {1{`RANDOM}};
  pipelineReg_tagValid_2_valid = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  pipelineReg_tagValid_3_tag = _RAND_6[19:0];
  _RAND_7 = {1{`RANDOM}};
  pipelineReg_tagValid_3_valid = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  pipelineReg_phyTag = _RAND_8[19:0];
  _RAND_9 = {1{`RANDOM}};
  pipelineReg_index = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  pipelineReg_bankIndex = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  pipelineReg_valid = _RAND_11[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      pipelineReg_tagValid_0_tag <= 20'h0;
    end else if (_T_1) begin
      pipelineReg_tagValid_0_tag <= io_in_tagValid_0_tag;
    end
    if (reset) begin
      pipelineReg_tagValid_0_valid <= 1'h0;
    end else if (_T_1) begin
      pipelineReg_tagValid_0_valid <= io_in_tagValid_0_valid;
    end
    if (reset) begin
      pipelineReg_tagValid_1_tag <= 20'h0;
    end else if (_T_1) begin
      pipelineReg_tagValid_1_tag <= io_in_tagValid_1_tag;
    end
    if (reset) begin
      pipelineReg_tagValid_1_valid <= 1'h0;
    end else if (_T_1) begin
      pipelineReg_tagValid_1_valid <= io_in_tagValid_1_valid;
    end
    if (reset) begin
      pipelineReg_tagValid_2_tag <= 20'h0;
    end else if (_T_1) begin
      pipelineReg_tagValid_2_tag <= io_in_tagValid_2_tag;
    end
    if (reset) begin
      pipelineReg_tagValid_2_valid <= 1'h0;
    end else if (_T_1) begin
      pipelineReg_tagValid_2_valid <= io_in_tagValid_2_valid;
    end
    if (reset) begin
      pipelineReg_tagValid_3_tag <= 20'h0;
    end else if (_T_1) begin
      pipelineReg_tagValid_3_tag <= io_in_tagValid_3_tag;
    end
    if (reset) begin
      pipelineReg_tagValid_3_valid <= 1'h0;
    end else if (_T_1) begin
      pipelineReg_tagValid_3_valid <= io_in_tagValid_3_valid;
    end
    if (reset) begin
      pipelineReg_phyTag <= 20'h0;
    end else if (_T_1) begin
      pipelineReg_phyTag <= io_in_phyTag;
    end
    if (reset) begin
      pipelineReg_index <= 8'h0;
    end else if (_T_1) begin
      pipelineReg_index <= io_in_index;
    end
    if (reset) begin
      pipelineReg_bankIndex <= 1'h0;
    end else if (_T_1) begin
      pipelineReg_bankIndex <= io_in_bankIndex;
    end
    if (reset) begin
      pipelineReg_valid <= 1'h0;
    end else if (_T_1) begin
      pipelineReg_valid <= io_in_valid;
    end
  end
endmodule
module MSHR(
  input         clock,
  input         reset,
  output        io_missAddr_ready,
  input         io_missAddr_valid,
  input  [19:0] io_missAddr_bits_tag,
  input  [7:0]  io_missAddr_bits_index,
  input         io_missAddr_bits_bankIndex,
  input         io_readyForWB,
  output        io_writeBack,
  output [19:0] io_mshrInfo_tag,
  output [7:0]  io_mshrInfo_index,
  output        io_mshrInfo_bankIndex
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [19:0] missEntryReg_tag; // @[MSHR.scala 31:29]
  reg [7:0] missEntryReg_index; // @[MSHR.scala 31:29]
  reg  missEntryReg_bankIndex; // @[MSHR.scala 31:29]
  reg  wbNext; // @[MSHR.scala 32:23]
  reg  state; // @[MSHR.scala 35:22]
  wire  _T_1 = ~state; // @[MSHR.scala 39:30]
  wire  _GEN_3 = io_missAddr_valid | state; // @[MSHR.scala 43:31]
  wire  _GEN_6 = state & io_readyForWB; // @[Conditional.scala 39:67]
  assign io_missAddr_ready = ~state; // @[MSHR.scala 39:21]
  assign io_writeBack = wbNext; // @[MSHR.scala 37:16]
  assign io_mshrInfo_tag = missEntryReg_tag; // @[MSHR.scala 38:15]
  assign io_mshrInfo_index = missEntryReg_index; // @[MSHR.scala 38:15]
  assign io_mshrInfo_bankIndex = missEntryReg_bankIndex; // @[MSHR.scala 38:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  missEntryReg_tag = _RAND_0[19:0];
  _RAND_1 = {1{`RANDOM}};
  missEntryReg_index = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  missEntryReg_bankIndex = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  wbNext = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  state = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      missEntryReg_tag <= 20'h0;
    end else if (_T_1) begin
      if (io_missAddr_valid) begin
        missEntryReg_tag <= io_missAddr_bits_tag;
      end
    end
    if (reset) begin
      missEntryReg_index <= 8'h0;
    end else if (_T_1) begin
      if (io_missAddr_valid) begin
        missEntryReg_index <= io_missAddr_bits_index;
      end
    end
    if (reset) begin
      missEntryReg_bankIndex <= 1'h0;
    end else if (_T_1) begin
      if (io_missAddr_valid) begin
        missEntryReg_bankIndex <= io_missAddr_bits_bankIndex;
      end
    end
    if (reset) begin
      wbNext <= 1'h0;
    end else if (_T_1) begin
      wbNext <= 1'h0;
    end else begin
      wbNext <= _GEN_6;
    end
    if (reset) begin
      state <= 1'h0;
    end else if (_T_1) begin
      state <= _GEN_3;
    end else if (state) begin
      if (io_readyForWB) begin
        state <= 1'h0;
      end
    end
  end
endmodule
module MissComparator(
  input  [19:0] io_tagValid_0_tag,
  input         io_tagValid_0_valid,
  input  [19:0] io_tagValid_1_tag,
  input         io_tagValid_1_valid,
  input  [19:0] io_tagValid_2_tag,
  input         io_tagValid_2_valid,
  input  [19:0] io_tagValid_3_tag,
  input         io_tagValid_3_valid,
  input  [19:0] io_phyTag,
  input  [7:0]  io_index,
  input  [19:0] io_mshr_bits_tag,
  input  [7:0]  io_mshr_bits_index,
  input         io_refillBufferValid,
  output        io_bankHitWay_valid,
  output [1:0]  io_bankHitWay_bits,
  output        io_hitInRefillBuffer
);
  wire  _T = io_tagValid_0_tag == io_phyTag; // @[MissComparator.scala 24:89]
  wire  bankHitVec_0 = io_tagValid_0_valid & _T; // @[MissComparator.scala 24:67]
  wire  _T_2 = io_tagValid_1_tag == io_phyTag; // @[MissComparator.scala 24:89]
  wire  bankHitVec_1 = io_tagValid_1_valid & _T_2; // @[MissComparator.scala 24:67]
  wire  _T_4 = io_tagValid_2_tag == io_phyTag; // @[MissComparator.scala 24:89]
  wire  bankHitVec_2 = io_tagValid_2_valid & _T_4; // @[MissComparator.scala 24:67]
  wire  _T_6 = io_tagValid_3_tag == io_phyTag; // @[MissComparator.scala 24:89]
  wire  bankHitVec_3 = io_tagValid_3_valid & _T_6; // @[MissComparator.scala 24:67]
  wire  _T_13 = bankHitVec_0 | bankHitVec_1; // @[MissComparator.scala 26:45]
  wire  _T_14 = _T_13 | bankHitVec_2; // @[MissComparator.scala 26:45]
  wire [1:0] _T_20 = bankHitVec_2 ? 2'h2 : 2'h3; // @[MissComparator.scala 27:46]
  wire [1:0] _T_21 = bankHitVec_1 ? 2'h1 : _T_20; // @[MissComparator.scala 27:46]
  wire  _T_23 = io_phyTag == io_mshr_bits_tag; // @[MissComparator.scala 34:15]
  wire  _T_24 = io_index == io_mshr_bits_index; // @[MissComparator.scala 35:16]
  wire  _T_25 = _T_23 & _T_24; // @[MissComparator.scala 34:36]
  assign io_bankHitWay_valid = _T_14 | bankHitVec_3; // @[MissComparator.scala 26:23]
  assign io_bankHitWay_bits = bankHitVec_0 ? 2'h0 : _T_21; // @[MissComparator.scala 27:22]
  assign io_hitInRefillBuffer = _T_25 & io_refillBufferValid; // @[MissComparator.scala 33:24]
endmodule
module AXIReadPort(
  input         clock,
  input         reset,
  input         io_axi_ar_ready,
  output        io_axi_ar_valid,
  output [31:0] io_axi_ar_bits_addr,
  output        io_axi_r_ready,
  input         io_axi_r_valid,
  input  [31:0] io_axi_r_bits_data,
  input         io_axi_r_bits_last,
  input         io_addrReq_valid,
  input  [31:0] io_addrReq_bits,
  output        io_transferData_valid,
  output [31:0] io_transferData_bits,
  output        io_finishTransfer
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] readState; // @[AXIReadPort.scala 30:26]
  wire  _T = readState == 2'h1; // @[AXIReadPort.scala 51:32]
  wire  _T_1 = readState == 2'h0; // @[AXIReadPort.scala 51:64]
  wire  _T_2 = _T_1 & io_addrReq_valid; // @[AXIReadPort.scala 51:77]
  wire  _T_4 = readState == 2'h2; // @[AXIReadPort.scala 52:31]
  wire  _T_6 = io_axi_r_ready & io_axi_r_valid; // @[Decoupled.scala 40:37]
  wire  _T_7 = _T_4 & _T_6; // @[AXIReadPort.scala 54:55]
  wire  _T_12 = 2'h0 == readState; // @[Conditional.scala 37:30]
  wire  _T_13 = io_axi_ar_ready & io_axi_ar_valid; // @[Decoupled.scala 40:37]
  wire  _T_15 = 2'h1 == readState; // @[Conditional.scala 37:30]
  wire  _T_17 = 2'h2 == readState; // @[Conditional.scala 37:30]
  wire  _T_19 = _T_6 & io_axi_r_bits_last; // @[AXIReadPort.scala 71:26]
  assign io_axi_ar_valid = _T | _T_2; // @[AXIReadPort.scala 51:19]
  assign io_axi_ar_bits_addr = io_addrReq_bits; // @[AXIReadPort.scala 37:23]
  assign io_axi_r_ready = readState == 2'h2; // @[AXIReadPort.scala 52:18]
  assign io_transferData_valid = _T_4 & _T_6; // @[AXIReadPort.scala 54:25]
  assign io_transferData_bits = io_axi_r_bits_data; // @[AXIReadPort.scala 55:24]
  assign io_finishTransfer = _T_7 & io_axi_r_bits_last; // @[AXIReadPort.scala 57:21]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  readState = _RAND_0[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      readState <= 2'h0;
    end else if (_T_12) begin
      if (io_addrReq_valid) begin
        if (_T_13) begin
          readState <= 2'h2;
        end else begin
          readState <= 2'h1;
        end
      end
    end else if (_T_15) begin
      if (_T_13) begin
        readState <= 2'h2;
      end
    end else if (_T_17) begin
      if (_T_19) begin
        readState <= 2'h0;
      end
    end
  end
endmodule
module ReFillBuffer(
  input         clock,
  input         reset,
  input         io_addr_valid,
  input         io_addr_bits,
  input         io_inputData_valid,
  input  [31:0] io_inputData_bits,
  input         io_finish,
  output        io_queryResult_valid,
  output [31:0] io_queryResult_bits,
  output [31:0] io_allData_0,
  output [31:0] io_allData_1
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  reg  state; // @[ReFillBuffer.scala 25:22]
  reg [31:0] buffer_0; // @[ReFillBuffer.scala 27:19]
  reg [31:0] buffer_1; // @[ReFillBuffer.scala 27:19]
  reg  bufferValidMask_0; // @[ReFillBuffer.scala 30:32]
  reg  bufferValidMask_1; // @[ReFillBuffer.scala 30:32]
  reg  writePtr; // @[ReFillBuffer.scala 32:21]
  wire  _T_1 = ~state; // @[Conditional.scala 37:30]
  wire  _GEN_7 = io_addr_valid | state; // @[ReFillBuffer.scala 41:27]
  wire  _T_6 = writePtr + 1'h1; // @[ReFillBuffer.scala 50:30]
  wire  _GEN_34 = ~writePtr; // @[ReFillBuffer.scala 51:35]
  wire  _GEN_10 = _GEN_34 | bufferValidMask_0; // @[ReFillBuffer.scala 51:35]
  wire  _GEN_11 = writePtr | bufferValidMask_1; // @[ReFillBuffer.scala 51:35]
  assign io_queryResult_valid = io_addr_bits ? bufferValidMask_1 : bufferValidMask_0; // @[ReFillBuffer.scala 34:24]
  assign io_queryResult_bits = io_addr_bits ? buffer_1 : buffer_0; // @[ReFillBuffer.scala 35:23]
  assign io_allData_0 = buffer_0; // @[ReFillBuffer.scala 37:14]
  assign io_allData_1 = buffer_1; // @[ReFillBuffer.scala 37:14]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  buffer_0 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  buffer_1 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  bufferValidMask_0 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  bufferValidMask_1 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  writePtr = _RAND_5[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      state <= 1'h0;
    end else if (_T_1) begin
      state <= _GEN_7;
    end else if (state) begin
      if (io_finish) begin
        state <= 1'h0;
      end
    end
    if (_T_1) begin
      if (io_addr_valid) begin
        buffer_0 <= 32'h0;
      end
    end else if (state) begin
      if (io_inputData_valid) begin
        if (~writePtr) begin
          buffer_0 <= io_inputData_bits;
        end
      end
    end
    if (_T_1) begin
      if (io_addr_valid) begin
        buffer_1 <= 32'h0;
      end
    end else if (state) begin
      if (io_inputData_valid) begin
        if (writePtr) begin
          buffer_1 <= io_inputData_bits;
        end
      end
    end
    if (reset) begin
      bufferValidMask_0 <= 1'h0;
    end else if (_T_1) begin
      if (io_addr_valid) begin
        bufferValidMask_0 <= 1'h0;
      end
    end else if (state) begin
      if (io_finish) begin
        bufferValidMask_0 <= 1'h0;
      end else if (io_inputData_valid) begin
        bufferValidMask_0 <= _GEN_10;
      end
    end
    if (reset) begin
      bufferValidMask_1 <= 1'h0;
    end else if (_T_1) begin
      if (io_addr_valid) begin
        bufferValidMask_1 <= 1'h0;
      end
    end else if (state) begin
      if (io_finish) begin
        bufferValidMask_1 <= 1'h0;
      end else if (io_inputData_valid) begin
        bufferValidMask_1 <= _GEN_11;
      end
    end
    if (_T_1) begin
      if (io_addr_valid) begin
        writePtr <= io_addr_bits;
      end
    end else if (state) begin
      if (io_inputData_valid) begin
        writePtr <= _T_6;
      end
    end
  end
endmodule
module ReadHolder(
  input         clock,
  input         reset,
  input         io_input_valid,
  input  [31:0] io_input_bits,
  output        io_output_valid,
  output [31:0] io_output_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] instruction; // @[ReadHolder.scala 16:28]
  reg  valid; // @[ReadHolder.scala 17:28]
  assign io_output_valid = valid; // @[ReadHolder.scala 22:19]
  assign io_output_bits = instruction; // @[ReadHolder.scala 20:19]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  instruction = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  valid = _RAND_1[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      instruction <= 32'h0;
    end else begin
      instruction <= io_input_bits;
    end
    if (reset) begin
      valid <= 1'h0;
    end else begin
      valid <= io_input_valid;
    end
  end
endmodule
module QueryTop(
  input         clock,
  input         reset,
  input         io_flush,
  output        io_ready,
  input  [19:0] io_fetchQuery_tagValid_0_tag,
  input         io_fetchQuery_tagValid_0_valid,
  input  [19:0] io_fetchQuery_tagValid_1_tag,
  input         io_fetchQuery_tagValid_1_valid,
  input  [19:0] io_fetchQuery_tagValid_2_tag,
  input         io_fetchQuery_tagValid_2_valid,
  input  [19:0] io_fetchQuery_tagValid_3_tag,
  input         io_fetchQuery_tagValid_3_valid,
  input  [19:0] io_fetchQuery_phyTag,
  input  [7:0]  io_fetchQuery_index,
  input         io_fetchQuery_bankIndex,
  input         io_fetchQuery_valid,
  input  [31:0] io_bankData_0,
  input  [31:0] io_bankData_1,
  input  [31:0] io_bankData_2,
  input  [31:0] io_bankData_3,
  input         io_data_ready,
  output        io_data_valid,
  output [31:0] io_data_bits,
  output        io_writeBundle_writeEnable,
  output [1:0]  io_writeBundle_writeWay,
  output [7:0]  io_writeBundle_writeIndex,
  output [19:0] io_writeBundle_writeTag,
  output [31:0] io_writeBundle_writeData_0,
  output [31:0] io_writeBundle_writeData_1,
  input         io_axi_ar_ready,
  output        io_axi_ar_valid,
  output [31:0] io_axi_ar_bits_addr,
  output        io_axi_r_ready,
  input         io_axi_r_valid,
  input  [31:0] io_axi_r_bits_data,
  input         io_axi_r_bits_last
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [31:0] _RAND_513;
  reg [31:0] _RAND_514;
  reg [31:0] _RAND_515;
  reg [31:0] _RAND_516;
  reg [31:0] _RAND_517;
  reg [31:0] _RAND_518;
  reg [31:0] _RAND_519;
  reg [31:0] _RAND_520;
  reg [31:0] _RAND_521;
  reg [31:0] _RAND_522;
  reg [31:0] _RAND_523;
  reg [31:0] _RAND_524;
  reg [31:0] _RAND_525;
  reg [31:0] _RAND_526;
  reg [31:0] _RAND_527;
  reg [31:0] _RAND_528;
  reg [31:0] _RAND_529;
  reg [31:0] _RAND_530;
  reg [31:0] _RAND_531;
  reg [31:0] _RAND_532;
  reg [31:0] _RAND_533;
  reg [31:0] _RAND_534;
  reg [31:0] _RAND_535;
  reg [31:0] _RAND_536;
  reg [31:0] _RAND_537;
  reg [31:0] _RAND_538;
  reg [31:0] _RAND_539;
  reg [31:0] _RAND_540;
  reg [31:0] _RAND_541;
  reg [31:0] _RAND_542;
  reg [31:0] _RAND_543;
  reg [31:0] _RAND_544;
  reg [31:0] _RAND_545;
  reg [31:0] _RAND_546;
  reg [31:0] _RAND_547;
  reg [31:0] _RAND_548;
  reg [31:0] _RAND_549;
  reg [31:0] _RAND_550;
  reg [31:0] _RAND_551;
  reg [31:0] _RAND_552;
  reg [31:0] _RAND_553;
  reg [31:0] _RAND_554;
  reg [31:0] _RAND_555;
  reg [31:0] _RAND_556;
  reg [31:0] _RAND_557;
  reg [31:0] _RAND_558;
  reg [31:0] _RAND_559;
  reg [31:0] _RAND_560;
  reg [31:0] _RAND_561;
  reg [31:0] _RAND_562;
  reg [31:0] _RAND_563;
  reg [31:0] _RAND_564;
  reg [31:0] _RAND_565;
  reg [31:0] _RAND_566;
  reg [31:0] _RAND_567;
  reg [31:0] _RAND_568;
  reg [31:0] _RAND_569;
  reg [31:0] _RAND_570;
  reg [31:0] _RAND_571;
  reg [31:0] _RAND_572;
  reg [31:0] _RAND_573;
  reg [31:0] _RAND_574;
  reg [31:0] _RAND_575;
  reg [31:0] _RAND_576;
  reg [31:0] _RAND_577;
  reg [31:0] _RAND_578;
  reg [31:0] _RAND_579;
  reg [31:0] _RAND_580;
  reg [31:0] _RAND_581;
  reg [31:0] _RAND_582;
  reg [31:0] _RAND_583;
  reg [31:0] _RAND_584;
  reg [31:0] _RAND_585;
  reg [31:0] _RAND_586;
  reg [31:0] _RAND_587;
  reg [31:0] _RAND_588;
  reg [31:0] _RAND_589;
  reg [31:0] _RAND_590;
  reg [31:0] _RAND_591;
  reg [31:0] _RAND_592;
  reg [31:0] _RAND_593;
  reg [31:0] _RAND_594;
  reg [31:0] _RAND_595;
  reg [31:0] _RAND_596;
  reg [31:0] _RAND_597;
  reg [31:0] _RAND_598;
  reg [31:0] _RAND_599;
  reg [31:0] _RAND_600;
  reg [31:0] _RAND_601;
  reg [31:0] _RAND_602;
  reg [31:0] _RAND_603;
  reg [31:0] _RAND_604;
  reg [31:0] _RAND_605;
  reg [31:0] _RAND_606;
  reg [31:0] _RAND_607;
  reg [31:0] _RAND_608;
  reg [31:0] _RAND_609;
  reg [31:0] _RAND_610;
  reg [31:0] _RAND_611;
  reg [31:0] _RAND_612;
  reg [31:0] _RAND_613;
  reg [31:0] _RAND_614;
  reg [31:0] _RAND_615;
  reg [31:0] _RAND_616;
  reg [31:0] _RAND_617;
  reg [31:0] _RAND_618;
  reg [31:0] _RAND_619;
  reg [31:0] _RAND_620;
  reg [31:0] _RAND_621;
  reg [31:0] _RAND_622;
  reg [31:0] _RAND_623;
  reg [31:0] _RAND_624;
  reg [31:0] _RAND_625;
  reg [31:0] _RAND_626;
  reg [31:0] _RAND_627;
  reg [31:0] _RAND_628;
  reg [31:0] _RAND_629;
  reg [31:0] _RAND_630;
  reg [31:0] _RAND_631;
  reg [31:0] _RAND_632;
  reg [31:0] _RAND_633;
  reg [31:0] _RAND_634;
  reg [31:0] _RAND_635;
  reg [31:0] _RAND_636;
  reg [31:0] _RAND_637;
  reg [31:0] _RAND_638;
  reg [31:0] _RAND_639;
  reg [31:0] _RAND_640;
  reg [31:0] _RAND_641;
  reg [31:0] _RAND_642;
  reg [31:0] _RAND_643;
  reg [31:0] _RAND_644;
  reg [31:0] _RAND_645;
  reg [31:0] _RAND_646;
  reg [31:0] _RAND_647;
  reg [31:0] _RAND_648;
  reg [31:0] _RAND_649;
  reg [31:0] _RAND_650;
  reg [31:0] _RAND_651;
  reg [31:0] _RAND_652;
  reg [31:0] _RAND_653;
  reg [31:0] _RAND_654;
  reg [31:0] _RAND_655;
  reg [31:0] _RAND_656;
  reg [31:0] _RAND_657;
  reg [31:0] _RAND_658;
  reg [31:0] _RAND_659;
  reg [31:0] _RAND_660;
  reg [31:0] _RAND_661;
  reg [31:0] _RAND_662;
  reg [31:0] _RAND_663;
  reg [31:0] _RAND_664;
  reg [31:0] _RAND_665;
  reg [31:0] _RAND_666;
  reg [31:0] _RAND_667;
  reg [31:0] _RAND_668;
  reg [31:0] _RAND_669;
  reg [31:0] _RAND_670;
  reg [31:0] _RAND_671;
  reg [31:0] _RAND_672;
  reg [31:0] _RAND_673;
  reg [31:0] _RAND_674;
  reg [31:0] _RAND_675;
  reg [31:0] _RAND_676;
  reg [31:0] _RAND_677;
  reg [31:0] _RAND_678;
  reg [31:0] _RAND_679;
  reg [31:0] _RAND_680;
  reg [31:0] _RAND_681;
  reg [31:0] _RAND_682;
  reg [31:0] _RAND_683;
  reg [31:0] _RAND_684;
  reg [31:0] _RAND_685;
  reg [31:0] _RAND_686;
  reg [31:0] _RAND_687;
  reg [31:0] _RAND_688;
  reg [31:0] _RAND_689;
  reg [31:0] _RAND_690;
  reg [31:0] _RAND_691;
  reg [31:0] _RAND_692;
  reg [31:0] _RAND_693;
  reg [31:0] _RAND_694;
  reg [31:0] _RAND_695;
  reg [31:0] _RAND_696;
  reg [31:0] _RAND_697;
  reg [31:0] _RAND_698;
  reg [31:0] _RAND_699;
  reg [31:0] _RAND_700;
  reg [31:0] _RAND_701;
  reg [31:0] _RAND_702;
  reg [31:0] _RAND_703;
  reg [31:0] _RAND_704;
  reg [31:0] _RAND_705;
  reg [31:0] _RAND_706;
  reg [31:0] _RAND_707;
  reg [31:0] _RAND_708;
  reg [31:0] _RAND_709;
  reg [31:0] _RAND_710;
  reg [31:0] _RAND_711;
  reg [31:0] _RAND_712;
  reg [31:0] _RAND_713;
  reg [31:0] _RAND_714;
  reg [31:0] _RAND_715;
  reg [31:0] _RAND_716;
  reg [31:0] _RAND_717;
  reg [31:0] _RAND_718;
  reg [31:0] _RAND_719;
  reg [31:0] _RAND_720;
  reg [31:0] _RAND_721;
  reg [31:0] _RAND_722;
  reg [31:0] _RAND_723;
  reg [31:0] _RAND_724;
  reg [31:0] _RAND_725;
  reg [31:0] _RAND_726;
  reg [31:0] _RAND_727;
  reg [31:0] _RAND_728;
  reg [31:0] _RAND_729;
  reg [31:0] _RAND_730;
  reg [31:0] _RAND_731;
  reg [31:0] _RAND_732;
  reg [31:0] _RAND_733;
  reg [31:0] _RAND_734;
  reg [31:0] _RAND_735;
  reg [31:0] _RAND_736;
  reg [31:0] _RAND_737;
  reg [31:0] _RAND_738;
  reg [31:0] _RAND_739;
  reg [31:0] _RAND_740;
  reg [31:0] _RAND_741;
  reg [31:0] _RAND_742;
  reg [31:0] _RAND_743;
  reg [31:0] _RAND_744;
  reg [31:0] _RAND_745;
  reg [31:0] _RAND_746;
  reg [31:0] _RAND_747;
  reg [31:0] _RAND_748;
  reg [31:0] _RAND_749;
  reg [31:0] _RAND_750;
  reg [31:0] _RAND_751;
  reg [31:0] _RAND_752;
  reg [31:0] _RAND_753;
  reg [31:0] _RAND_754;
  reg [31:0] _RAND_755;
  reg [31:0] _RAND_756;
  reg [31:0] _RAND_757;
  reg [31:0] _RAND_758;
  reg [31:0] _RAND_759;
  reg [31:0] _RAND_760;
  reg [31:0] _RAND_761;
  reg [31:0] _RAND_762;
  reg [31:0] _RAND_763;
  reg [31:0] _RAND_764;
  reg [31:0] _RAND_765;
  reg [31:0] _RAND_766;
  reg [31:0] _RAND_767;
  reg [31:0] _RAND_768;
  reg [31:0] _RAND_769;
  reg [31:0] _RAND_770;
  reg [31:0] _RAND_771;
  reg [31:0] _RAND_772;
  reg [31:0] _RAND_773;
  reg [31:0] _RAND_774;
  reg [31:0] _RAND_775;
  reg [31:0] _RAND_776;
  reg [31:0] _RAND_777;
  reg [31:0] _RAND_778;
  reg [31:0] _RAND_779;
  reg [31:0] _RAND_780;
  reg [31:0] _RAND_781;
  reg [31:0] _RAND_782;
  reg [31:0] _RAND_783;
  reg [31:0] _RAND_784;
  reg [31:0] _RAND_785;
  reg [31:0] _RAND_786;
  reg [31:0] _RAND_787;
  reg [31:0] _RAND_788;
  reg [31:0] _RAND_789;
  reg [31:0] _RAND_790;
  reg [31:0] _RAND_791;
  reg [31:0] _RAND_792;
  reg [31:0] _RAND_793;
  reg [31:0] _RAND_794;
  reg [31:0] _RAND_795;
  reg [31:0] _RAND_796;
  reg [31:0] _RAND_797;
  reg [31:0] _RAND_798;
  reg [31:0] _RAND_799;
  reg [31:0] _RAND_800;
  reg [31:0] _RAND_801;
  reg [31:0] _RAND_802;
  reg [31:0] _RAND_803;
  reg [31:0] _RAND_804;
  reg [31:0] _RAND_805;
  reg [31:0] _RAND_806;
  reg [31:0] _RAND_807;
  reg [31:0] _RAND_808;
  reg [31:0] _RAND_809;
  reg [31:0] _RAND_810;
  reg [31:0] _RAND_811;
  reg [31:0] _RAND_812;
  reg [31:0] _RAND_813;
  reg [31:0] _RAND_814;
  reg [31:0] _RAND_815;
  reg [31:0] _RAND_816;
  reg [31:0] _RAND_817;
  reg [31:0] _RAND_818;
  reg [31:0] _RAND_819;
  reg [31:0] _RAND_820;
  reg [31:0] _RAND_821;
  reg [31:0] _RAND_822;
  reg [31:0] _RAND_823;
  reg [31:0] _RAND_824;
  reg [31:0] _RAND_825;
  reg [31:0] _RAND_826;
  reg [31:0] _RAND_827;
  reg [31:0] _RAND_828;
  reg [31:0] _RAND_829;
  reg [31:0] _RAND_830;
  reg [31:0] _RAND_831;
  reg [31:0] _RAND_832;
  reg [31:0] _RAND_833;
  reg [31:0] _RAND_834;
  reg [31:0] _RAND_835;
  reg [31:0] _RAND_836;
  reg [31:0] _RAND_837;
  reg [31:0] _RAND_838;
  reg [31:0] _RAND_839;
  reg [31:0] _RAND_840;
  reg [31:0] _RAND_841;
  reg [31:0] _RAND_842;
  reg [31:0] _RAND_843;
  reg [31:0] _RAND_844;
  reg [31:0] _RAND_845;
  reg [31:0] _RAND_846;
  reg [31:0] _RAND_847;
  reg [31:0] _RAND_848;
  reg [31:0] _RAND_849;
  reg [31:0] _RAND_850;
  reg [31:0] _RAND_851;
  reg [31:0] _RAND_852;
  reg [31:0] _RAND_853;
  reg [31:0] _RAND_854;
  reg [31:0] _RAND_855;
  reg [31:0] _RAND_856;
  reg [31:0] _RAND_857;
  reg [31:0] _RAND_858;
  reg [31:0] _RAND_859;
  reg [31:0] _RAND_860;
  reg [31:0] _RAND_861;
  reg [31:0] _RAND_862;
  reg [31:0] _RAND_863;
  reg [31:0] _RAND_864;
  reg [31:0] _RAND_865;
  reg [31:0] _RAND_866;
  reg [31:0] _RAND_867;
  reg [31:0] _RAND_868;
  reg [31:0] _RAND_869;
  reg [31:0] _RAND_870;
  reg [31:0] _RAND_871;
  reg [31:0] _RAND_872;
  reg [31:0] _RAND_873;
  reg [31:0] _RAND_874;
  reg [31:0] _RAND_875;
  reg [31:0] _RAND_876;
  reg [31:0] _RAND_877;
  reg [31:0] _RAND_878;
  reg [31:0] _RAND_879;
  reg [31:0] _RAND_880;
  reg [31:0] _RAND_881;
  reg [31:0] _RAND_882;
  reg [31:0] _RAND_883;
  reg [31:0] _RAND_884;
  reg [31:0] _RAND_885;
  reg [31:0] _RAND_886;
  reg [31:0] _RAND_887;
  reg [31:0] _RAND_888;
  reg [31:0] _RAND_889;
  reg [31:0] _RAND_890;
  reg [31:0] _RAND_891;
  reg [31:0] _RAND_892;
  reg [31:0] _RAND_893;
  reg [31:0] _RAND_894;
  reg [31:0] _RAND_895;
  reg [31:0] _RAND_896;
  reg [31:0] _RAND_897;
  reg [31:0] _RAND_898;
  reg [31:0] _RAND_899;
  reg [31:0] _RAND_900;
  reg [31:0] _RAND_901;
  reg [31:0] _RAND_902;
  reg [31:0] _RAND_903;
  reg [31:0] _RAND_904;
  reg [31:0] _RAND_905;
  reg [31:0] _RAND_906;
  reg [31:0] _RAND_907;
  reg [31:0] _RAND_908;
  reg [31:0] _RAND_909;
  reg [31:0] _RAND_910;
  reg [31:0] _RAND_911;
  reg [31:0] _RAND_912;
  reg [31:0] _RAND_913;
  reg [31:0] _RAND_914;
  reg [31:0] _RAND_915;
  reg [31:0] _RAND_916;
  reg [31:0] _RAND_917;
  reg [31:0] _RAND_918;
  reg [31:0] _RAND_919;
  reg [31:0] _RAND_920;
  reg [31:0] _RAND_921;
  reg [31:0] _RAND_922;
  reg [31:0] _RAND_923;
  reg [31:0] _RAND_924;
  reg [31:0] _RAND_925;
  reg [31:0] _RAND_926;
  reg [31:0] _RAND_927;
  reg [31:0] _RAND_928;
  reg [31:0] _RAND_929;
  reg [31:0] _RAND_930;
  reg [31:0] _RAND_931;
  reg [31:0] _RAND_932;
  reg [31:0] _RAND_933;
  reg [31:0] _RAND_934;
  reg [31:0] _RAND_935;
  reg [31:0] _RAND_936;
  reg [31:0] _RAND_937;
  reg [31:0] _RAND_938;
  reg [31:0] _RAND_939;
  reg [31:0] _RAND_940;
  reg [31:0] _RAND_941;
  reg [31:0] _RAND_942;
  reg [31:0] _RAND_943;
  reg [31:0] _RAND_944;
  reg [31:0] _RAND_945;
  reg [31:0] _RAND_946;
  reg [31:0] _RAND_947;
  reg [31:0] _RAND_948;
  reg [31:0] _RAND_949;
  reg [31:0] _RAND_950;
  reg [31:0] _RAND_951;
  reg [31:0] _RAND_952;
  reg [31:0] _RAND_953;
  reg [31:0] _RAND_954;
  reg [31:0] _RAND_955;
  reg [31:0] _RAND_956;
  reg [31:0] _RAND_957;
  reg [31:0] _RAND_958;
  reg [31:0] _RAND_959;
  reg [31:0] _RAND_960;
  reg [31:0] _RAND_961;
  reg [31:0] _RAND_962;
  reg [31:0] _RAND_963;
  reg [31:0] _RAND_964;
  reg [31:0] _RAND_965;
  reg [31:0] _RAND_966;
  reg [31:0] _RAND_967;
  reg [31:0] _RAND_968;
  reg [31:0] _RAND_969;
  reg [31:0] _RAND_970;
  reg [31:0] _RAND_971;
  reg [31:0] _RAND_972;
  reg [31:0] _RAND_973;
  reg [31:0] _RAND_974;
  reg [31:0] _RAND_975;
  reg [31:0] _RAND_976;
  reg [31:0] _RAND_977;
  reg [31:0] _RAND_978;
  reg [31:0] _RAND_979;
  reg [31:0] _RAND_980;
  reg [31:0] _RAND_981;
  reg [31:0] _RAND_982;
  reg [31:0] _RAND_983;
  reg [31:0] _RAND_984;
  reg [31:0] _RAND_985;
  reg [31:0] _RAND_986;
  reg [31:0] _RAND_987;
  reg [31:0] _RAND_988;
  reg [31:0] _RAND_989;
  reg [31:0] _RAND_990;
  reg [31:0] _RAND_991;
  reg [31:0] _RAND_992;
  reg [31:0] _RAND_993;
  reg [31:0] _RAND_994;
  reg [31:0] _RAND_995;
  reg [31:0] _RAND_996;
  reg [31:0] _RAND_997;
  reg [31:0] _RAND_998;
  reg [31:0] _RAND_999;
  reg [31:0] _RAND_1000;
  reg [31:0] _RAND_1001;
  reg [31:0] _RAND_1002;
  reg [31:0] _RAND_1003;
  reg [31:0] _RAND_1004;
  reg [31:0] _RAND_1005;
  reg [31:0] _RAND_1006;
  reg [31:0] _RAND_1007;
  reg [31:0] _RAND_1008;
  reg [31:0] _RAND_1009;
  reg [31:0] _RAND_1010;
  reg [31:0] _RAND_1011;
  reg [31:0] _RAND_1012;
  reg [31:0] _RAND_1013;
  reg [31:0] _RAND_1014;
  reg [31:0] _RAND_1015;
  reg [31:0] _RAND_1016;
  reg [31:0] _RAND_1017;
  reg [31:0] _RAND_1018;
  reg [31:0] _RAND_1019;
  reg [31:0] _RAND_1020;
  reg [31:0] _RAND_1021;
  reg [31:0] _RAND_1022;
  reg [31:0] _RAND_1023;
`endif // RANDOMIZE_REG_INIT
  wire  mshr_clock; // @[QueryTop.scala 37:28]
  wire  mshr_reset; // @[QueryTop.scala 37:28]
  wire  mshr_io_missAddr_ready; // @[QueryTop.scala 37:28]
  wire  mshr_io_missAddr_valid; // @[QueryTop.scala 37:28]
  wire [19:0] mshr_io_missAddr_bits_tag; // @[QueryTop.scala 37:28]
  wire [7:0] mshr_io_missAddr_bits_index; // @[QueryTop.scala 37:28]
  wire  mshr_io_missAddr_bits_bankIndex; // @[QueryTop.scala 37:28]
  wire  mshr_io_readyForWB; // @[QueryTop.scala 37:28]
  wire  mshr_io_writeBack; // @[QueryTop.scala 37:28]
  wire [19:0] mshr_io_mshrInfo_tag; // @[QueryTop.scala 37:28]
  wire [7:0] mshr_io_mshrInfo_index; // @[QueryTop.scala 37:28]
  wire  mshr_io_mshrInfo_bankIndex; // @[QueryTop.scala 37:28]
  wire [19:0] comparator_io_tagValid_0_tag; // @[QueryTop.scala 38:28]
  wire  comparator_io_tagValid_0_valid; // @[QueryTop.scala 38:28]
  wire [19:0] comparator_io_tagValid_1_tag; // @[QueryTop.scala 38:28]
  wire  comparator_io_tagValid_1_valid; // @[QueryTop.scala 38:28]
  wire [19:0] comparator_io_tagValid_2_tag; // @[QueryTop.scala 38:28]
  wire  comparator_io_tagValid_2_valid; // @[QueryTop.scala 38:28]
  wire [19:0] comparator_io_tagValid_3_tag; // @[QueryTop.scala 38:28]
  wire  comparator_io_tagValid_3_valid; // @[QueryTop.scala 38:28]
  wire [19:0] comparator_io_phyTag; // @[QueryTop.scala 38:28]
  wire [7:0] comparator_io_index; // @[QueryTop.scala 38:28]
  wire [19:0] comparator_io_mshr_bits_tag; // @[QueryTop.scala 38:28]
  wire [7:0] comparator_io_mshr_bits_index; // @[QueryTop.scala 38:28]
  wire  comparator_io_refillBufferValid; // @[QueryTop.scala 38:28]
  wire  comparator_io_bankHitWay_valid; // @[QueryTop.scala 38:28]
  wire [1:0] comparator_io_bankHitWay_bits; // @[QueryTop.scala 38:28]
  wire  comparator_io_hitInRefillBuffer; // @[QueryTop.scala 38:28]
  wire  axi_clock; // @[QueryTop.scala 39:28]
  wire  axi_reset; // @[QueryTop.scala 39:28]
  wire  axi_io_axi_ar_ready; // @[QueryTop.scala 39:28]
  wire  axi_io_axi_ar_valid; // @[QueryTop.scala 39:28]
  wire [31:0] axi_io_axi_ar_bits_addr; // @[QueryTop.scala 39:28]
  wire  axi_io_axi_r_ready; // @[QueryTop.scala 39:28]
  wire  axi_io_axi_r_valid; // @[QueryTop.scala 39:28]
  wire [31:0] axi_io_axi_r_bits_data; // @[QueryTop.scala 39:28]
  wire  axi_io_axi_r_bits_last; // @[QueryTop.scala 39:28]
  wire  axi_io_addrReq_valid; // @[QueryTop.scala 39:28]
  wire [31:0] axi_io_addrReq_bits; // @[QueryTop.scala 39:28]
  wire  axi_io_transferData_valid; // @[QueryTop.scala 39:28]
  wire [31:0] axi_io_transferData_bits; // @[QueryTop.scala 39:28]
  wire  axi_io_finishTransfer; // @[QueryTop.scala 39:28]
  wire  refillBuffer_clock; // @[QueryTop.scala 40:28]
  wire  refillBuffer_reset; // @[QueryTop.scala 40:28]
  wire  refillBuffer_io_addr_valid; // @[QueryTop.scala 40:28]
  wire  refillBuffer_io_addr_bits; // @[QueryTop.scala 40:28]
  wire  refillBuffer_io_inputData_valid; // @[QueryTop.scala 40:28]
  wire [31:0] refillBuffer_io_inputData_bits; // @[QueryTop.scala 40:28]
  wire  refillBuffer_io_finish; // @[QueryTop.scala 40:28]
  wire  refillBuffer_io_queryResult_valid; // @[QueryTop.scala 40:28]
  wire [31:0] refillBuffer_io_queryResult_bits; // @[QueryTop.scala 40:28]
  wire [31:0] refillBuffer_io_allData_0; // @[QueryTop.scala 40:28]
  wire [31:0] refillBuffer_io_allData_1; // @[QueryTop.scala 40:28]
  wire  readHolder_clock; // @[QueryTop.scala 42:28]
  wire  readHolder_reset; // @[QueryTop.scala 42:28]
  wire  readHolder_io_input_valid; // @[QueryTop.scala 42:28]
  wire [31:0] readHolder_io_input_bits; // @[QueryTop.scala 42:28]
  wire  readHolder_io_output_valid; // @[QueryTop.scala 42:28]
  wire [31:0] readHolder_io_output_bits; // @[QueryTop.scala 42:28]
  reg  _T_257_0_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_0_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_0_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_0_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_1_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_1_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_1_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_1_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_2_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_2_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_2_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_2_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_3_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_3_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_3_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_3_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_4_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_4_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_4_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_4_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_5_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_5_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_5_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_5_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_6_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_6_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_6_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_6_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_7_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_7_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_7_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_7_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_8_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_8_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_8_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_8_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_9_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_9_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_9_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_9_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_10_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_10_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_10_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_10_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_11_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_11_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_11_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_11_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_12_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_12_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_12_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_12_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_13_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_13_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_13_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_13_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_14_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_14_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_14_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_14_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_15_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_15_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_15_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_15_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_16_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_16_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_16_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_16_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_17_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_17_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_17_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_17_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_18_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_18_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_18_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_18_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_19_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_19_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_19_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_19_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_20_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_20_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_20_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_20_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_21_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_21_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_21_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_21_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_22_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_22_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_22_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_22_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_23_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_23_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_23_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_23_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_24_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_24_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_24_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_24_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_25_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_25_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_25_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_25_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_26_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_26_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_26_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_26_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_27_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_27_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_27_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_27_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_28_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_28_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_28_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_28_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_29_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_29_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_29_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_29_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_30_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_30_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_30_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_30_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_31_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_31_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_31_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_31_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_32_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_32_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_32_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_32_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_33_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_33_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_33_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_33_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_34_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_34_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_34_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_34_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_35_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_35_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_35_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_35_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_36_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_36_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_36_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_36_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_37_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_37_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_37_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_37_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_38_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_38_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_38_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_38_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_39_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_39_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_39_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_39_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_40_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_40_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_40_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_40_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_41_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_41_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_41_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_41_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_42_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_42_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_42_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_42_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_43_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_43_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_43_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_43_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_44_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_44_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_44_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_44_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_45_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_45_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_45_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_45_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_46_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_46_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_46_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_46_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_47_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_47_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_47_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_47_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_48_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_48_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_48_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_48_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_49_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_49_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_49_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_49_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_50_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_50_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_50_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_50_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_51_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_51_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_51_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_51_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_52_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_52_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_52_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_52_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_53_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_53_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_53_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_53_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_54_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_54_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_54_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_54_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_55_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_55_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_55_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_55_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_56_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_56_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_56_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_56_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_57_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_57_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_57_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_57_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_58_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_58_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_58_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_58_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_59_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_59_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_59_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_59_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_60_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_60_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_60_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_60_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_61_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_61_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_61_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_61_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_62_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_62_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_62_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_62_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_63_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_63_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_63_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_63_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_64_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_64_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_64_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_64_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_65_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_65_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_65_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_65_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_66_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_66_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_66_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_66_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_67_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_67_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_67_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_67_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_68_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_68_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_68_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_68_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_69_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_69_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_69_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_69_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_70_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_70_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_70_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_70_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_71_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_71_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_71_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_71_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_72_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_72_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_72_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_72_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_73_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_73_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_73_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_73_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_74_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_74_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_74_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_74_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_75_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_75_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_75_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_75_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_76_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_76_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_76_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_76_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_77_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_77_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_77_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_77_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_78_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_78_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_78_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_78_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_79_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_79_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_79_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_79_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_80_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_80_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_80_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_80_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_81_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_81_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_81_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_81_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_82_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_82_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_82_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_82_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_83_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_83_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_83_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_83_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_84_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_84_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_84_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_84_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_85_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_85_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_85_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_85_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_86_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_86_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_86_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_86_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_87_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_87_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_87_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_87_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_88_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_88_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_88_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_88_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_89_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_89_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_89_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_89_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_90_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_90_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_90_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_90_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_91_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_91_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_91_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_91_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_92_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_92_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_92_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_92_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_93_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_93_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_93_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_93_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_94_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_94_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_94_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_94_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_95_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_95_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_95_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_95_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_96_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_96_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_96_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_96_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_97_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_97_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_97_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_97_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_98_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_98_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_98_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_98_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_99_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_99_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_99_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_99_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_100_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_100_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_100_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_100_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_101_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_101_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_101_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_101_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_102_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_102_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_102_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_102_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_103_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_103_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_103_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_103_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_104_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_104_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_104_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_104_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_105_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_105_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_105_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_105_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_106_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_106_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_106_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_106_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_107_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_107_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_107_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_107_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_108_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_108_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_108_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_108_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_109_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_109_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_109_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_109_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_110_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_110_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_110_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_110_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_111_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_111_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_111_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_111_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_112_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_112_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_112_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_112_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_113_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_113_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_113_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_113_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_114_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_114_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_114_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_114_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_115_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_115_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_115_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_115_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_116_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_116_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_116_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_116_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_117_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_117_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_117_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_117_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_118_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_118_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_118_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_118_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_119_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_119_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_119_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_119_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_120_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_120_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_120_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_120_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_121_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_121_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_121_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_121_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_122_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_122_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_122_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_122_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_123_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_123_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_123_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_123_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_124_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_124_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_124_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_124_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_125_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_125_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_125_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_125_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_126_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_126_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_126_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_126_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_127_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_127_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_127_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_127_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_128_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_128_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_128_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_128_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_129_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_129_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_129_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_129_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_130_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_130_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_130_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_130_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_131_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_131_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_131_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_131_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_132_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_132_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_132_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_132_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_133_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_133_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_133_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_133_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_134_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_134_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_134_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_134_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_135_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_135_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_135_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_135_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_136_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_136_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_136_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_136_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_137_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_137_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_137_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_137_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_138_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_138_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_138_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_138_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_139_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_139_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_139_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_139_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_140_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_140_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_140_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_140_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_141_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_141_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_141_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_141_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_142_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_142_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_142_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_142_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_143_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_143_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_143_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_143_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_144_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_144_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_144_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_144_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_145_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_145_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_145_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_145_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_146_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_146_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_146_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_146_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_147_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_147_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_147_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_147_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_148_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_148_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_148_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_148_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_149_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_149_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_149_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_149_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_150_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_150_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_150_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_150_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_151_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_151_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_151_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_151_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_152_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_152_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_152_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_152_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_153_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_153_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_153_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_153_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_154_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_154_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_154_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_154_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_155_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_155_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_155_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_155_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_156_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_156_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_156_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_156_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_157_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_157_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_157_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_157_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_158_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_158_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_158_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_158_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_159_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_159_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_159_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_159_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_160_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_160_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_160_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_160_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_161_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_161_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_161_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_161_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_162_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_162_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_162_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_162_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_163_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_163_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_163_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_163_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_164_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_164_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_164_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_164_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_165_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_165_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_165_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_165_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_166_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_166_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_166_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_166_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_167_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_167_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_167_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_167_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_168_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_168_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_168_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_168_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_169_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_169_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_169_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_169_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_170_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_170_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_170_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_170_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_171_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_171_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_171_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_171_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_172_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_172_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_172_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_172_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_173_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_173_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_173_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_173_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_174_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_174_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_174_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_174_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_175_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_175_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_175_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_175_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_176_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_176_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_176_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_176_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_177_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_177_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_177_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_177_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_178_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_178_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_178_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_178_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_179_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_179_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_179_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_179_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_180_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_180_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_180_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_180_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_181_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_181_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_181_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_181_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_182_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_182_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_182_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_182_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_183_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_183_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_183_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_183_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_184_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_184_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_184_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_184_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_185_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_185_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_185_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_185_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_186_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_186_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_186_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_186_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_187_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_187_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_187_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_187_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_188_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_188_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_188_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_188_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_189_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_189_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_189_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_189_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_190_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_190_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_190_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_190_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_191_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_191_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_191_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_191_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_192_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_192_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_192_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_192_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_193_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_193_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_193_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_193_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_194_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_194_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_194_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_194_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_195_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_195_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_195_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_195_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_196_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_196_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_196_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_196_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_197_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_197_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_197_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_197_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_198_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_198_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_198_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_198_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_199_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_199_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_199_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_199_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_200_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_200_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_200_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_200_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_201_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_201_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_201_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_201_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_202_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_202_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_202_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_202_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_203_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_203_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_203_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_203_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_204_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_204_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_204_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_204_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_205_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_205_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_205_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_205_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_206_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_206_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_206_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_206_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_207_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_207_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_207_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_207_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_208_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_208_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_208_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_208_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_209_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_209_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_209_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_209_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_210_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_210_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_210_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_210_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_211_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_211_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_211_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_211_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_212_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_212_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_212_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_212_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_213_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_213_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_213_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_213_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_214_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_214_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_214_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_214_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_215_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_215_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_215_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_215_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_216_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_216_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_216_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_216_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_217_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_217_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_217_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_217_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_218_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_218_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_218_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_218_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_219_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_219_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_219_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_219_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_220_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_220_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_220_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_220_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_221_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_221_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_221_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_221_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_222_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_222_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_222_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_222_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_223_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_223_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_223_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_223_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_224_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_224_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_224_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_224_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_225_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_225_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_225_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_225_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_226_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_226_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_226_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_226_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_227_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_227_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_227_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_227_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_228_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_228_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_228_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_228_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_229_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_229_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_229_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_229_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_230_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_230_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_230_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_230_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_231_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_231_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_231_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_231_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_232_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_232_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_232_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_232_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_233_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_233_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_233_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_233_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_234_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_234_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_234_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_234_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_235_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_235_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_235_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_235_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_236_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_236_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_236_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_236_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_237_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_237_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_237_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_237_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_238_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_238_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_238_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_238_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_239_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_239_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_239_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_239_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_240_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_240_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_240_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_240_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_241_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_241_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_241_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_241_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_242_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_242_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_242_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_242_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_243_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_243_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_243_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_243_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_244_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_244_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_244_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_244_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_245_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_245_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_245_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_245_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_246_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_246_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_246_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_246_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_247_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_247_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_247_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_247_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_248_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_248_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_248_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_248_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_249_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_249_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_249_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_249_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_250_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_250_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_250_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_250_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_251_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_251_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_251_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_251_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_252_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_252_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_252_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_252_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_253_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_253_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_253_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_253_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_254_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_254_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_254_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_254_3; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_255_0; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_255_1; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_255_2; // @[PLRUMRUNM.scala 15:23]
  reg  _T_257_255_3; // @[PLRUMRUNM.scala 15:23]
  wire  _T_258 = ~io_fetchQuery_valid; // @[QueryTop.scala 45:33]
  wire  passThrough = _T_258 | io_flush; // @[QueryTop.scala 45:54]
  wire  newMiss = mshr_io_missAddr_ready & mshr_io_missAddr_valid; // @[Decoupled.scala 40:37]
  wire  hitInBank = comparator_io_bankHitWay_valid;
  wire  hitInRefillBuffer = comparator_io_hitInRefillBuffer;
  wire  queryHit = hitInBank | hitInRefillBuffer; // @[QueryTop.scala 57:40]
  wire  _T_262 = ~passThrough; // @[QueryTop.scala 60:43]
  wire  validData = queryHit & _T_262; // @[QueryTop.scala 60:40]
  wire  _T_264 = io_data_ready & io_data_valid; // @[Decoupled.scala 40:37]
  wire [31:0] _GEN_1 = 2'h1 == comparator_io_bankHitWay_bits ? io_bankData_1 : io_bankData_0; // @[Mux.scala 98:16]
  wire [31:0] _GEN_2 = 2'h2 == comparator_io_bankHitWay_bits ? io_bankData_2 : _GEN_1; // @[Mux.scala 98:16]
  wire [31:0] _GEN_3 = 2'h3 == comparator_io_bankHitWay_bits ? io_bankData_3 : _GEN_2; // @[Mux.scala 98:16]
  wire [31:0] _T_266 = comparator_io_hitInRefillBuffer ? refillBuffer_io_queryResult_bits : _GEN_3; // @[Mux.scala 98:16]
  wire  _GEN_9 = 8'h1 == mshr_io_mshrInfo_index ? _T_257_1_1 : _T_257_0_1;
  wire  _GEN_10 = 8'h1 == mshr_io_mshrInfo_index ? _T_257_1_2 : _T_257_0_2;
  wire  _GEN_11 = 8'h1 == mshr_io_mshrInfo_index ? _T_257_1_3 : _T_257_0_3;
  wire  _GEN_13 = 8'h2 == mshr_io_mshrInfo_index ? _T_257_2_1 : _GEN_9;
  wire  _GEN_14 = 8'h2 == mshr_io_mshrInfo_index ? _T_257_2_2 : _GEN_10;
  wire  _GEN_15 = 8'h2 == mshr_io_mshrInfo_index ? _T_257_2_3 : _GEN_11;
  wire  _GEN_17 = 8'h3 == mshr_io_mshrInfo_index ? _T_257_3_1 : _GEN_13;
  wire  _GEN_18 = 8'h3 == mshr_io_mshrInfo_index ? _T_257_3_2 : _GEN_14;
  wire  _GEN_19 = 8'h3 == mshr_io_mshrInfo_index ? _T_257_3_3 : _GEN_15;
  wire  _GEN_21 = 8'h4 == mshr_io_mshrInfo_index ? _T_257_4_1 : _GEN_17;
  wire  _GEN_22 = 8'h4 == mshr_io_mshrInfo_index ? _T_257_4_2 : _GEN_18;
  wire  _GEN_23 = 8'h4 == mshr_io_mshrInfo_index ? _T_257_4_3 : _GEN_19;
  wire  _GEN_25 = 8'h5 == mshr_io_mshrInfo_index ? _T_257_5_1 : _GEN_21;
  wire  _GEN_26 = 8'h5 == mshr_io_mshrInfo_index ? _T_257_5_2 : _GEN_22;
  wire  _GEN_27 = 8'h5 == mshr_io_mshrInfo_index ? _T_257_5_3 : _GEN_23;
  wire  _GEN_29 = 8'h6 == mshr_io_mshrInfo_index ? _T_257_6_1 : _GEN_25;
  wire  _GEN_30 = 8'h6 == mshr_io_mshrInfo_index ? _T_257_6_2 : _GEN_26;
  wire  _GEN_31 = 8'h6 == mshr_io_mshrInfo_index ? _T_257_6_3 : _GEN_27;
  wire  _GEN_33 = 8'h7 == mshr_io_mshrInfo_index ? _T_257_7_1 : _GEN_29;
  wire  _GEN_34 = 8'h7 == mshr_io_mshrInfo_index ? _T_257_7_2 : _GEN_30;
  wire  _GEN_35 = 8'h7 == mshr_io_mshrInfo_index ? _T_257_7_3 : _GEN_31;
  wire  _GEN_37 = 8'h8 == mshr_io_mshrInfo_index ? _T_257_8_1 : _GEN_33;
  wire  _GEN_38 = 8'h8 == mshr_io_mshrInfo_index ? _T_257_8_2 : _GEN_34;
  wire  _GEN_39 = 8'h8 == mshr_io_mshrInfo_index ? _T_257_8_3 : _GEN_35;
  wire  _GEN_41 = 8'h9 == mshr_io_mshrInfo_index ? _T_257_9_1 : _GEN_37;
  wire  _GEN_42 = 8'h9 == mshr_io_mshrInfo_index ? _T_257_9_2 : _GEN_38;
  wire  _GEN_43 = 8'h9 == mshr_io_mshrInfo_index ? _T_257_9_3 : _GEN_39;
  wire  _GEN_45 = 8'ha == mshr_io_mshrInfo_index ? _T_257_10_1 : _GEN_41;
  wire  _GEN_46 = 8'ha == mshr_io_mshrInfo_index ? _T_257_10_2 : _GEN_42;
  wire  _GEN_47 = 8'ha == mshr_io_mshrInfo_index ? _T_257_10_3 : _GEN_43;
  wire  _GEN_49 = 8'hb == mshr_io_mshrInfo_index ? _T_257_11_1 : _GEN_45;
  wire  _GEN_50 = 8'hb == mshr_io_mshrInfo_index ? _T_257_11_2 : _GEN_46;
  wire  _GEN_51 = 8'hb == mshr_io_mshrInfo_index ? _T_257_11_3 : _GEN_47;
  wire  _GEN_53 = 8'hc == mshr_io_mshrInfo_index ? _T_257_12_1 : _GEN_49;
  wire  _GEN_54 = 8'hc == mshr_io_mshrInfo_index ? _T_257_12_2 : _GEN_50;
  wire  _GEN_55 = 8'hc == mshr_io_mshrInfo_index ? _T_257_12_3 : _GEN_51;
  wire  _GEN_57 = 8'hd == mshr_io_mshrInfo_index ? _T_257_13_1 : _GEN_53;
  wire  _GEN_58 = 8'hd == mshr_io_mshrInfo_index ? _T_257_13_2 : _GEN_54;
  wire  _GEN_59 = 8'hd == mshr_io_mshrInfo_index ? _T_257_13_3 : _GEN_55;
  wire  _GEN_61 = 8'he == mshr_io_mshrInfo_index ? _T_257_14_1 : _GEN_57;
  wire  _GEN_62 = 8'he == mshr_io_mshrInfo_index ? _T_257_14_2 : _GEN_58;
  wire  _GEN_63 = 8'he == mshr_io_mshrInfo_index ? _T_257_14_3 : _GEN_59;
  wire  _GEN_65 = 8'hf == mshr_io_mshrInfo_index ? _T_257_15_1 : _GEN_61;
  wire  _GEN_66 = 8'hf == mshr_io_mshrInfo_index ? _T_257_15_2 : _GEN_62;
  wire  _GEN_67 = 8'hf == mshr_io_mshrInfo_index ? _T_257_15_3 : _GEN_63;
  wire  _GEN_69 = 8'h10 == mshr_io_mshrInfo_index ? _T_257_16_1 : _GEN_65;
  wire  _GEN_70 = 8'h10 == mshr_io_mshrInfo_index ? _T_257_16_2 : _GEN_66;
  wire  _GEN_71 = 8'h10 == mshr_io_mshrInfo_index ? _T_257_16_3 : _GEN_67;
  wire  _GEN_73 = 8'h11 == mshr_io_mshrInfo_index ? _T_257_17_1 : _GEN_69;
  wire  _GEN_74 = 8'h11 == mshr_io_mshrInfo_index ? _T_257_17_2 : _GEN_70;
  wire  _GEN_75 = 8'h11 == mshr_io_mshrInfo_index ? _T_257_17_3 : _GEN_71;
  wire  _GEN_77 = 8'h12 == mshr_io_mshrInfo_index ? _T_257_18_1 : _GEN_73;
  wire  _GEN_78 = 8'h12 == mshr_io_mshrInfo_index ? _T_257_18_2 : _GEN_74;
  wire  _GEN_79 = 8'h12 == mshr_io_mshrInfo_index ? _T_257_18_3 : _GEN_75;
  wire  _GEN_81 = 8'h13 == mshr_io_mshrInfo_index ? _T_257_19_1 : _GEN_77;
  wire  _GEN_82 = 8'h13 == mshr_io_mshrInfo_index ? _T_257_19_2 : _GEN_78;
  wire  _GEN_83 = 8'h13 == mshr_io_mshrInfo_index ? _T_257_19_3 : _GEN_79;
  wire  _GEN_85 = 8'h14 == mshr_io_mshrInfo_index ? _T_257_20_1 : _GEN_81;
  wire  _GEN_86 = 8'h14 == mshr_io_mshrInfo_index ? _T_257_20_2 : _GEN_82;
  wire  _GEN_87 = 8'h14 == mshr_io_mshrInfo_index ? _T_257_20_3 : _GEN_83;
  wire  _GEN_89 = 8'h15 == mshr_io_mshrInfo_index ? _T_257_21_1 : _GEN_85;
  wire  _GEN_90 = 8'h15 == mshr_io_mshrInfo_index ? _T_257_21_2 : _GEN_86;
  wire  _GEN_91 = 8'h15 == mshr_io_mshrInfo_index ? _T_257_21_3 : _GEN_87;
  wire  _GEN_93 = 8'h16 == mshr_io_mshrInfo_index ? _T_257_22_1 : _GEN_89;
  wire  _GEN_94 = 8'h16 == mshr_io_mshrInfo_index ? _T_257_22_2 : _GEN_90;
  wire  _GEN_95 = 8'h16 == mshr_io_mshrInfo_index ? _T_257_22_3 : _GEN_91;
  wire  _GEN_97 = 8'h17 == mshr_io_mshrInfo_index ? _T_257_23_1 : _GEN_93;
  wire  _GEN_98 = 8'h17 == mshr_io_mshrInfo_index ? _T_257_23_2 : _GEN_94;
  wire  _GEN_99 = 8'h17 == mshr_io_mshrInfo_index ? _T_257_23_3 : _GEN_95;
  wire  _GEN_101 = 8'h18 == mshr_io_mshrInfo_index ? _T_257_24_1 : _GEN_97;
  wire  _GEN_102 = 8'h18 == mshr_io_mshrInfo_index ? _T_257_24_2 : _GEN_98;
  wire  _GEN_103 = 8'h18 == mshr_io_mshrInfo_index ? _T_257_24_3 : _GEN_99;
  wire  _GEN_105 = 8'h19 == mshr_io_mshrInfo_index ? _T_257_25_1 : _GEN_101;
  wire  _GEN_106 = 8'h19 == mshr_io_mshrInfo_index ? _T_257_25_2 : _GEN_102;
  wire  _GEN_107 = 8'h19 == mshr_io_mshrInfo_index ? _T_257_25_3 : _GEN_103;
  wire  _GEN_109 = 8'h1a == mshr_io_mshrInfo_index ? _T_257_26_1 : _GEN_105;
  wire  _GEN_110 = 8'h1a == mshr_io_mshrInfo_index ? _T_257_26_2 : _GEN_106;
  wire  _GEN_111 = 8'h1a == mshr_io_mshrInfo_index ? _T_257_26_3 : _GEN_107;
  wire  _GEN_113 = 8'h1b == mshr_io_mshrInfo_index ? _T_257_27_1 : _GEN_109;
  wire  _GEN_114 = 8'h1b == mshr_io_mshrInfo_index ? _T_257_27_2 : _GEN_110;
  wire  _GEN_115 = 8'h1b == mshr_io_mshrInfo_index ? _T_257_27_3 : _GEN_111;
  wire  _GEN_117 = 8'h1c == mshr_io_mshrInfo_index ? _T_257_28_1 : _GEN_113;
  wire  _GEN_118 = 8'h1c == mshr_io_mshrInfo_index ? _T_257_28_2 : _GEN_114;
  wire  _GEN_119 = 8'h1c == mshr_io_mshrInfo_index ? _T_257_28_3 : _GEN_115;
  wire  _GEN_121 = 8'h1d == mshr_io_mshrInfo_index ? _T_257_29_1 : _GEN_117;
  wire  _GEN_122 = 8'h1d == mshr_io_mshrInfo_index ? _T_257_29_2 : _GEN_118;
  wire  _GEN_123 = 8'h1d == mshr_io_mshrInfo_index ? _T_257_29_3 : _GEN_119;
  wire  _GEN_125 = 8'h1e == mshr_io_mshrInfo_index ? _T_257_30_1 : _GEN_121;
  wire  _GEN_126 = 8'h1e == mshr_io_mshrInfo_index ? _T_257_30_2 : _GEN_122;
  wire  _GEN_127 = 8'h1e == mshr_io_mshrInfo_index ? _T_257_30_3 : _GEN_123;
  wire  _GEN_129 = 8'h1f == mshr_io_mshrInfo_index ? _T_257_31_1 : _GEN_125;
  wire  _GEN_130 = 8'h1f == mshr_io_mshrInfo_index ? _T_257_31_2 : _GEN_126;
  wire  _GEN_131 = 8'h1f == mshr_io_mshrInfo_index ? _T_257_31_3 : _GEN_127;
  wire  _GEN_133 = 8'h20 == mshr_io_mshrInfo_index ? _T_257_32_1 : _GEN_129;
  wire  _GEN_134 = 8'h20 == mshr_io_mshrInfo_index ? _T_257_32_2 : _GEN_130;
  wire  _GEN_135 = 8'h20 == mshr_io_mshrInfo_index ? _T_257_32_3 : _GEN_131;
  wire  _GEN_137 = 8'h21 == mshr_io_mshrInfo_index ? _T_257_33_1 : _GEN_133;
  wire  _GEN_138 = 8'h21 == mshr_io_mshrInfo_index ? _T_257_33_2 : _GEN_134;
  wire  _GEN_139 = 8'h21 == mshr_io_mshrInfo_index ? _T_257_33_3 : _GEN_135;
  wire  _GEN_141 = 8'h22 == mshr_io_mshrInfo_index ? _T_257_34_1 : _GEN_137;
  wire  _GEN_142 = 8'h22 == mshr_io_mshrInfo_index ? _T_257_34_2 : _GEN_138;
  wire  _GEN_143 = 8'h22 == mshr_io_mshrInfo_index ? _T_257_34_3 : _GEN_139;
  wire  _GEN_145 = 8'h23 == mshr_io_mshrInfo_index ? _T_257_35_1 : _GEN_141;
  wire  _GEN_146 = 8'h23 == mshr_io_mshrInfo_index ? _T_257_35_2 : _GEN_142;
  wire  _GEN_147 = 8'h23 == mshr_io_mshrInfo_index ? _T_257_35_3 : _GEN_143;
  wire  _GEN_149 = 8'h24 == mshr_io_mshrInfo_index ? _T_257_36_1 : _GEN_145;
  wire  _GEN_150 = 8'h24 == mshr_io_mshrInfo_index ? _T_257_36_2 : _GEN_146;
  wire  _GEN_151 = 8'h24 == mshr_io_mshrInfo_index ? _T_257_36_3 : _GEN_147;
  wire  _GEN_153 = 8'h25 == mshr_io_mshrInfo_index ? _T_257_37_1 : _GEN_149;
  wire  _GEN_154 = 8'h25 == mshr_io_mshrInfo_index ? _T_257_37_2 : _GEN_150;
  wire  _GEN_155 = 8'h25 == mshr_io_mshrInfo_index ? _T_257_37_3 : _GEN_151;
  wire  _GEN_157 = 8'h26 == mshr_io_mshrInfo_index ? _T_257_38_1 : _GEN_153;
  wire  _GEN_158 = 8'h26 == mshr_io_mshrInfo_index ? _T_257_38_2 : _GEN_154;
  wire  _GEN_159 = 8'h26 == mshr_io_mshrInfo_index ? _T_257_38_3 : _GEN_155;
  wire  _GEN_161 = 8'h27 == mshr_io_mshrInfo_index ? _T_257_39_1 : _GEN_157;
  wire  _GEN_162 = 8'h27 == mshr_io_mshrInfo_index ? _T_257_39_2 : _GEN_158;
  wire  _GEN_163 = 8'h27 == mshr_io_mshrInfo_index ? _T_257_39_3 : _GEN_159;
  wire  _GEN_165 = 8'h28 == mshr_io_mshrInfo_index ? _T_257_40_1 : _GEN_161;
  wire  _GEN_166 = 8'h28 == mshr_io_mshrInfo_index ? _T_257_40_2 : _GEN_162;
  wire  _GEN_167 = 8'h28 == mshr_io_mshrInfo_index ? _T_257_40_3 : _GEN_163;
  wire  _GEN_169 = 8'h29 == mshr_io_mshrInfo_index ? _T_257_41_1 : _GEN_165;
  wire  _GEN_170 = 8'h29 == mshr_io_mshrInfo_index ? _T_257_41_2 : _GEN_166;
  wire  _GEN_171 = 8'h29 == mshr_io_mshrInfo_index ? _T_257_41_3 : _GEN_167;
  wire  _GEN_173 = 8'h2a == mshr_io_mshrInfo_index ? _T_257_42_1 : _GEN_169;
  wire  _GEN_174 = 8'h2a == mshr_io_mshrInfo_index ? _T_257_42_2 : _GEN_170;
  wire  _GEN_175 = 8'h2a == mshr_io_mshrInfo_index ? _T_257_42_3 : _GEN_171;
  wire  _GEN_177 = 8'h2b == mshr_io_mshrInfo_index ? _T_257_43_1 : _GEN_173;
  wire  _GEN_178 = 8'h2b == mshr_io_mshrInfo_index ? _T_257_43_2 : _GEN_174;
  wire  _GEN_179 = 8'h2b == mshr_io_mshrInfo_index ? _T_257_43_3 : _GEN_175;
  wire  _GEN_181 = 8'h2c == mshr_io_mshrInfo_index ? _T_257_44_1 : _GEN_177;
  wire  _GEN_182 = 8'h2c == mshr_io_mshrInfo_index ? _T_257_44_2 : _GEN_178;
  wire  _GEN_183 = 8'h2c == mshr_io_mshrInfo_index ? _T_257_44_3 : _GEN_179;
  wire  _GEN_185 = 8'h2d == mshr_io_mshrInfo_index ? _T_257_45_1 : _GEN_181;
  wire  _GEN_186 = 8'h2d == mshr_io_mshrInfo_index ? _T_257_45_2 : _GEN_182;
  wire  _GEN_187 = 8'h2d == mshr_io_mshrInfo_index ? _T_257_45_3 : _GEN_183;
  wire  _GEN_189 = 8'h2e == mshr_io_mshrInfo_index ? _T_257_46_1 : _GEN_185;
  wire  _GEN_190 = 8'h2e == mshr_io_mshrInfo_index ? _T_257_46_2 : _GEN_186;
  wire  _GEN_191 = 8'h2e == mshr_io_mshrInfo_index ? _T_257_46_3 : _GEN_187;
  wire  _GEN_193 = 8'h2f == mshr_io_mshrInfo_index ? _T_257_47_1 : _GEN_189;
  wire  _GEN_194 = 8'h2f == mshr_io_mshrInfo_index ? _T_257_47_2 : _GEN_190;
  wire  _GEN_195 = 8'h2f == mshr_io_mshrInfo_index ? _T_257_47_3 : _GEN_191;
  wire  _GEN_197 = 8'h30 == mshr_io_mshrInfo_index ? _T_257_48_1 : _GEN_193;
  wire  _GEN_198 = 8'h30 == mshr_io_mshrInfo_index ? _T_257_48_2 : _GEN_194;
  wire  _GEN_199 = 8'h30 == mshr_io_mshrInfo_index ? _T_257_48_3 : _GEN_195;
  wire  _GEN_201 = 8'h31 == mshr_io_mshrInfo_index ? _T_257_49_1 : _GEN_197;
  wire  _GEN_202 = 8'h31 == mshr_io_mshrInfo_index ? _T_257_49_2 : _GEN_198;
  wire  _GEN_203 = 8'h31 == mshr_io_mshrInfo_index ? _T_257_49_3 : _GEN_199;
  wire  _GEN_205 = 8'h32 == mshr_io_mshrInfo_index ? _T_257_50_1 : _GEN_201;
  wire  _GEN_206 = 8'h32 == mshr_io_mshrInfo_index ? _T_257_50_2 : _GEN_202;
  wire  _GEN_207 = 8'h32 == mshr_io_mshrInfo_index ? _T_257_50_3 : _GEN_203;
  wire  _GEN_209 = 8'h33 == mshr_io_mshrInfo_index ? _T_257_51_1 : _GEN_205;
  wire  _GEN_210 = 8'h33 == mshr_io_mshrInfo_index ? _T_257_51_2 : _GEN_206;
  wire  _GEN_211 = 8'h33 == mshr_io_mshrInfo_index ? _T_257_51_3 : _GEN_207;
  wire  _GEN_213 = 8'h34 == mshr_io_mshrInfo_index ? _T_257_52_1 : _GEN_209;
  wire  _GEN_214 = 8'h34 == mshr_io_mshrInfo_index ? _T_257_52_2 : _GEN_210;
  wire  _GEN_215 = 8'h34 == mshr_io_mshrInfo_index ? _T_257_52_3 : _GEN_211;
  wire  _GEN_217 = 8'h35 == mshr_io_mshrInfo_index ? _T_257_53_1 : _GEN_213;
  wire  _GEN_218 = 8'h35 == mshr_io_mshrInfo_index ? _T_257_53_2 : _GEN_214;
  wire  _GEN_219 = 8'h35 == mshr_io_mshrInfo_index ? _T_257_53_3 : _GEN_215;
  wire  _GEN_221 = 8'h36 == mshr_io_mshrInfo_index ? _T_257_54_1 : _GEN_217;
  wire  _GEN_222 = 8'h36 == mshr_io_mshrInfo_index ? _T_257_54_2 : _GEN_218;
  wire  _GEN_223 = 8'h36 == mshr_io_mshrInfo_index ? _T_257_54_3 : _GEN_219;
  wire  _GEN_225 = 8'h37 == mshr_io_mshrInfo_index ? _T_257_55_1 : _GEN_221;
  wire  _GEN_226 = 8'h37 == mshr_io_mshrInfo_index ? _T_257_55_2 : _GEN_222;
  wire  _GEN_227 = 8'h37 == mshr_io_mshrInfo_index ? _T_257_55_3 : _GEN_223;
  wire  _GEN_229 = 8'h38 == mshr_io_mshrInfo_index ? _T_257_56_1 : _GEN_225;
  wire  _GEN_230 = 8'h38 == mshr_io_mshrInfo_index ? _T_257_56_2 : _GEN_226;
  wire  _GEN_231 = 8'h38 == mshr_io_mshrInfo_index ? _T_257_56_3 : _GEN_227;
  wire  _GEN_233 = 8'h39 == mshr_io_mshrInfo_index ? _T_257_57_1 : _GEN_229;
  wire  _GEN_234 = 8'h39 == mshr_io_mshrInfo_index ? _T_257_57_2 : _GEN_230;
  wire  _GEN_235 = 8'h39 == mshr_io_mshrInfo_index ? _T_257_57_3 : _GEN_231;
  wire  _GEN_237 = 8'h3a == mshr_io_mshrInfo_index ? _T_257_58_1 : _GEN_233;
  wire  _GEN_238 = 8'h3a == mshr_io_mshrInfo_index ? _T_257_58_2 : _GEN_234;
  wire  _GEN_239 = 8'h3a == mshr_io_mshrInfo_index ? _T_257_58_3 : _GEN_235;
  wire  _GEN_241 = 8'h3b == mshr_io_mshrInfo_index ? _T_257_59_1 : _GEN_237;
  wire  _GEN_242 = 8'h3b == mshr_io_mshrInfo_index ? _T_257_59_2 : _GEN_238;
  wire  _GEN_243 = 8'h3b == mshr_io_mshrInfo_index ? _T_257_59_3 : _GEN_239;
  wire  _GEN_245 = 8'h3c == mshr_io_mshrInfo_index ? _T_257_60_1 : _GEN_241;
  wire  _GEN_246 = 8'h3c == mshr_io_mshrInfo_index ? _T_257_60_2 : _GEN_242;
  wire  _GEN_247 = 8'h3c == mshr_io_mshrInfo_index ? _T_257_60_3 : _GEN_243;
  wire  _GEN_249 = 8'h3d == mshr_io_mshrInfo_index ? _T_257_61_1 : _GEN_245;
  wire  _GEN_250 = 8'h3d == mshr_io_mshrInfo_index ? _T_257_61_2 : _GEN_246;
  wire  _GEN_251 = 8'h3d == mshr_io_mshrInfo_index ? _T_257_61_3 : _GEN_247;
  wire  _GEN_253 = 8'h3e == mshr_io_mshrInfo_index ? _T_257_62_1 : _GEN_249;
  wire  _GEN_254 = 8'h3e == mshr_io_mshrInfo_index ? _T_257_62_2 : _GEN_250;
  wire  _GEN_255 = 8'h3e == mshr_io_mshrInfo_index ? _T_257_62_3 : _GEN_251;
  wire  _GEN_257 = 8'h3f == mshr_io_mshrInfo_index ? _T_257_63_1 : _GEN_253;
  wire  _GEN_258 = 8'h3f == mshr_io_mshrInfo_index ? _T_257_63_2 : _GEN_254;
  wire  _GEN_259 = 8'h3f == mshr_io_mshrInfo_index ? _T_257_63_3 : _GEN_255;
  wire  _GEN_261 = 8'h40 == mshr_io_mshrInfo_index ? _T_257_64_1 : _GEN_257;
  wire  _GEN_262 = 8'h40 == mshr_io_mshrInfo_index ? _T_257_64_2 : _GEN_258;
  wire  _GEN_263 = 8'h40 == mshr_io_mshrInfo_index ? _T_257_64_3 : _GEN_259;
  wire  _GEN_265 = 8'h41 == mshr_io_mshrInfo_index ? _T_257_65_1 : _GEN_261;
  wire  _GEN_266 = 8'h41 == mshr_io_mshrInfo_index ? _T_257_65_2 : _GEN_262;
  wire  _GEN_267 = 8'h41 == mshr_io_mshrInfo_index ? _T_257_65_3 : _GEN_263;
  wire  _GEN_269 = 8'h42 == mshr_io_mshrInfo_index ? _T_257_66_1 : _GEN_265;
  wire  _GEN_270 = 8'h42 == mshr_io_mshrInfo_index ? _T_257_66_2 : _GEN_266;
  wire  _GEN_271 = 8'h42 == mshr_io_mshrInfo_index ? _T_257_66_3 : _GEN_267;
  wire  _GEN_273 = 8'h43 == mshr_io_mshrInfo_index ? _T_257_67_1 : _GEN_269;
  wire  _GEN_274 = 8'h43 == mshr_io_mshrInfo_index ? _T_257_67_2 : _GEN_270;
  wire  _GEN_275 = 8'h43 == mshr_io_mshrInfo_index ? _T_257_67_3 : _GEN_271;
  wire  _GEN_277 = 8'h44 == mshr_io_mshrInfo_index ? _T_257_68_1 : _GEN_273;
  wire  _GEN_278 = 8'h44 == mshr_io_mshrInfo_index ? _T_257_68_2 : _GEN_274;
  wire  _GEN_279 = 8'h44 == mshr_io_mshrInfo_index ? _T_257_68_3 : _GEN_275;
  wire  _GEN_281 = 8'h45 == mshr_io_mshrInfo_index ? _T_257_69_1 : _GEN_277;
  wire  _GEN_282 = 8'h45 == mshr_io_mshrInfo_index ? _T_257_69_2 : _GEN_278;
  wire  _GEN_283 = 8'h45 == mshr_io_mshrInfo_index ? _T_257_69_3 : _GEN_279;
  wire  _GEN_285 = 8'h46 == mshr_io_mshrInfo_index ? _T_257_70_1 : _GEN_281;
  wire  _GEN_286 = 8'h46 == mshr_io_mshrInfo_index ? _T_257_70_2 : _GEN_282;
  wire  _GEN_287 = 8'h46 == mshr_io_mshrInfo_index ? _T_257_70_3 : _GEN_283;
  wire  _GEN_289 = 8'h47 == mshr_io_mshrInfo_index ? _T_257_71_1 : _GEN_285;
  wire  _GEN_290 = 8'h47 == mshr_io_mshrInfo_index ? _T_257_71_2 : _GEN_286;
  wire  _GEN_291 = 8'h47 == mshr_io_mshrInfo_index ? _T_257_71_3 : _GEN_287;
  wire  _GEN_293 = 8'h48 == mshr_io_mshrInfo_index ? _T_257_72_1 : _GEN_289;
  wire  _GEN_294 = 8'h48 == mshr_io_mshrInfo_index ? _T_257_72_2 : _GEN_290;
  wire  _GEN_295 = 8'h48 == mshr_io_mshrInfo_index ? _T_257_72_3 : _GEN_291;
  wire  _GEN_297 = 8'h49 == mshr_io_mshrInfo_index ? _T_257_73_1 : _GEN_293;
  wire  _GEN_298 = 8'h49 == mshr_io_mshrInfo_index ? _T_257_73_2 : _GEN_294;
  wire  _GEN_299 = 8'h49 == mshr_io_mshrInfo_index ? _T_257_73_3 : _GEN_295;
  wire  _GEN_301 = 8'h4a == mshr_io_mshrInfo_index ? _T_257_74_1 : _GEN_297;
  wire  _GEN_302 = 8'h4a == mshr_io_mshrInfo_index ? _T_257_74_2 : _GEN_298;
  wire  _GEN_303 = 8'h4a == mshr_io_mshrInfo_index ? _T_257_74_3 : _GEN_299;
  wire  _GEN_305 = 8'h4b == mshr_io_mshrInfo_index ? _T_257_75_1 : _GEN_301;
  wire  _GEN_306 = 8'h4b == mshr_io_mshrInfo_index ? _T_257_75_2 : _GEN_302;
  wire  _GEN_307 = 8'h4b == mshr_io_mshrInfo_index ? _T_257_75_3 : _GEN_303;
  wire  _GEN_309 = 8'h4c == mshr_io_mshrInfo_index ? _T_257_76_1 : _GEN_305;
  wire  _GEN_310 = 8'h4c == mshr_io_mshrInfo_index ? _T_257_76_2 : _GEN_306;
  wire  _GEN_311 = 8'h4c == mshr_io_mshrInfo_index ? _T_257_76_3 : _GEN_307;
  wire  _GEN_313 = 8'h4d == mshr_io_mshrInfo_index ? _T_257_77_1 : _GEN_309;
  wire  _GEN_314 = 8'h4d == mshr_io_mshrInfo_index ? _T_257_77_2 : _GEN_310;
  wire  _GEN_315 = 8'h4d == mshr_io_mshrInfo_index ? _T_257_77_3 : _GEN_311;
  wire  _GEN_317 = 8'h4e == mshr_io_mshrInfo_index ? _T_257_78_1 : _GEN_313;
  wire  _GEN_318 = 8'h4e == mshr_io_mshrInfo_index ? _T_257_78_2 : _GEN_314;
  wire  _GEN_319 = 8'h4e == mshr_io_mshrInfo_index ? _T_257_78_3 : _GEN_315;
  wire  _GEN_321 = 8'h4f == mshr_io_mshrInfo_index ? _T_257_79_1 : _GEN_317;
  wire  _GEN_322 = 8'h4f == mshr_io_mshrInfo_index ? _T_257_79_2 : _GEN_318;
  wire  _GEN_323 = 8'h4f == mshr_io_mshrInfo_index ? _T_257_79_3 : _GEN_319;
  wire  _GEN_325 = 8'h50 == mshr_io_mshrInfo_index ? _T_257_80_1 : _GEN_321;
  wire  _GEN_326 = 8'h50 == mshr_io_mshrInfo_index ? _T_257_80_2 : _GEN_322;
  wire  _GEN_327 = 8'h50 == mshr_io_mshrInfo_index ? _T_257_80_3 : _GEN_323;
  wire  _GEN_329 = 8'h51 == mshr_io_mshrInfo_index ? _T_257_81_1 : _GEN_325;
  wire  _GEN_330 = 8'h51 == mshr_io_mshrInfo_index ? _T_257_81_2 : _GEN_326;
  wire  _GEN_331 = 8'h51 == mshr_io_mshrInfo_index ? _T_257_81_3 : _GEN_327;
  wire  _GEN_333 = 8'h52 == mshr_io_mshrInfo_index ? _T_257_82_1 : _GEN_329;
  wire  _GEN_334 = 8'h52 == mshr_io_mshrInfo_index ? _T_257_82_2 : _GEN_330;
  wire  _GEN_335 = 8'h52 == mshr_io_mshrInfo_index ? _T_257_82_3 : _GEN_331;
  wire  _GEN_337 = 8'h53 == mshr_io_mshrInfo_index ? _T_257_83_1 : _GEN_333;
  wire  _GEN_338 = 8'h53 == mshr_io_mshrInfo_index ? _T_257_83_2 : _GEN_334;
  wire  _GEN_339 = 8'h53 == mshr_io_mshrInfo_index ? _T_257_83_3 : _GEN_335;
  wire  _GEN_341 = 8'h54 == mshr_io_mshrInfo_index ? _T_257_84_1 : _GEN_337;
  wire  _GEN_342 = 8'h54 == mshr_io_mshrInfo_index ? _T_257_84_2 : _GEN_338;
  wire  _GEN_343 = 8'h54 == mshr_io_mshrInfo_index ? _T_257_84_3 : _GEN_339;
  wire  _GEN_345 = 8'h55 == mshr_io_mshrInfo_index ? _T_257_85_1 : _GEN_341;
  wire  _GEN_346 = 8'h55 == mshr_io_mshrInfo_index ? _T_257_85_2 : _GEN_342;
  wire  _GEN_347 = 8'h55 == mshr_io_mshrInfo_index ? _T_257_85_3 : _GEN_343;
  wire  _GEN_349 = 8'h56 == mshr_io_mshrInfo_index ? _T_257_86_1 : _GEN_345;
  wire  _GEN_350 = 8'h56 == mshr_io_mshrInfo_index ? _T_257_86_2 : _GEN_346;
  wire  _GEN_351 = 8'h56 == mshr_io_mshrInfo_index ? _T_257_86_3 : _GEN_347;
  wire  _GEN_353 = 8'h57 == mshr_io_mshrInfo_index ? _T_257_87_1 : _GEN_349;
  wire  _GEN_354 = 8'h57 == mshr_io_mshrInfo_index ? _T_257_87_2 : _GEN_350;
  wire  _GEN_355 = 8'h57 == mshr_io_mshrInfo_index ? _T_257_87_3 : _GEN_351;
  wire  _GEN_357 = 8'h58 == mshr_io_mshrInfo_index ? _T_257_88_1 : _GEN_353;
  wire  _GEN_358 = 8'h58 == mshr_io_mshrInfo_index ? _T_257_88_2 : _GEN_354;
  wire  _GEN_359 = 8'h58 == mshr_io_mshrInfo_index ? _T_257_88_3 : _GEN_355;
  wire  _GEN_361 = 8'h59 == mshr_io_mshrInfo_index ? _T_257_89_1 : _GEN_357;
  wire  _GEN_362 = 8'h59 == mshr_io_mshrInfo_index ? _T_257_89_2 : _GEN_358;
  wire  _GEN_363 = 8'h59 == mshr_io_mshrInfo_index ? _T_257_89_3 : _GEN_359;
  wire  _GEN_365 = 8'h5a == mshr_io_mshrInfo_index ? _T_257_90_1 : _GEN_361;
  wire  _GEN_366 = 8'h5a == mshr_io_mshrInfo_index ? _T_257_90_2 : _GEN_362;
  wire  _GEN_367 = 8'h5a == mshr_io_mshrInfo_index ? _T_257_90_3 : _GEN_363;
  wire  _GEN_369 = 8'h5b == mshr_io_mshrInfo_index ? _T_257_91_1 : _GEN_365;
  wire  _GEN_370 = 8'h5b == mshr_io_mshrInfo_index ? _T_257_91_2 : _GEN_366;
  wire  _GEN_371 = 8'h5b == mshr_io_mshrInfo_index ? _T_257_91_3 : _GEN_367;
  wire  _GEN_373 = 8'h5c == mshr_io_mshrInfo_index ? _T_257_92_1 : _GEN_369;
  wire  _GEN_374 = 8'h5c == mshr_io_mshrInfo_index ? _T_257_92_2 : _GEN_370;
  wire  _GEN_375 = 8'h5c == mshr_io_mshrInfo_index ? _T_257_92_3 : _GEN_371;
  wire  _GEN_377 = 8'h5d == mshr_io_mshrInfo_index ? _T_257_93_1 : _GEN_373;
  wire  _GEN_378 = 8'h5d == mshr_io_mshrInfo_index ? _T_257_93_2 : _GEN_374;
  wire  _GEN_379 = 8'h5d == mshr_io_mshrInfo_index ? _T_257_93_3 : _GEN_375;
  wire  _GEN_381 = 8'h5e == mshr_io_mshrInfo_index ? _T_257_94_1 : _GEN_377;
  wire  _GEN_382 = 8'h5e == mshr_io_mshrInfo_index ? _T_257_94_2 : _GEN_378;
  wire  _GEN_383 = 8'h5e == mshr_io_mshrInfo_index ? _T_257_94_3 : _GEN_379;
  wire  _GEN_385 = 8'h5f == mshr_io_mshrInfo_index ? _T_257_95_1 : _GEN_381;
  wire  _GEN_386 = 8'h5f == mshr_io_mshrInfo_index ? _T_257_95_2 : _GEN_382;
  wire  _GEN_387 = 8'h5f == mshr_io_mshrInfo_index ? _T_257_95_3 : _GEN_383;
  wire  _GEN_389 = 8'h60 == mshr_io_mshrInfo_index ? _T_257_96_1 : _GEN_385;
  wire  _GEN_390 = 8'h60 == mshr_io_mshrInfo_index ? _T_257_96_2 : _GEN_386;
  wire  _GEN_391 = 8'h60 == mshr_io_mshrInfo_index ? _T_257_96_3 : _GEN_387;
  wire  _GEN_393 = 8'h61 == mshr_io_mshrInfo_index ? _T_257_97_1 : _GEN_389;
  wire  _GEN_394 = 8'h61 == mshr_io_mshrInfo_index ? _T_257_97_2 : _GEN_390;
  wire  _GEN_395 = 8'h61 == mshr_io_mshrInfo_index ? _T_257_97_3 : _GEN_391;
  wire  _GEN_397 = 8'h62 == mshr_io_mshrInfo_index ? _T_257_98_1 : _GEN_393;
  wire  _GEN_398 = 8'h62 == mshr_io_mshrInfo_index ? _T_257_98_2 : _GEN_394;
  wire  _GEN_399 = 8'h62 == mshr_io_mshrInfo_index ? _T_257_98_3 : _GEN_395;
  wire  _GEN_401 = 8'h63 == mshr_io_mshrInfo_index ? _T_257_99_1 : _GEN_397;
  wire  _GEN_402 = 8'h63 == mshr_io_mshrInfo_index ? _T_257_99_2 : _GEN_398;
  wire  _GEN_403 = 8'h63 == mshr_io_mshrInfo_index ? _T_257_99_3 : _GEN_399;
  wire  _GEN_405 = 8'h64 == mshr_io_mshrInfo_index ? _T_257_100_1 : _GEN_401;
  wire  _GEN_406 = 8'h64 == mshr_io_mshrInfo_index ? _T_257_100_2 : _GEN_402;
  wire  _GEN_407 = 8'h64 == mshr_io_mshrInfo_index ? _T_257_100_3 : _GEN_403;
  wire  _GEN_409 = 8'h65 == mshr_io_mshrInfo_index ? _T_257_101_1 : _GEN_405;
  wire  _GEN_410 = 8'h65 == mshr_io_mshrInfo_index ? _T_257_101_2 : _GEN_406;
  wire  _GEN_411 = 8'h65 == mshr_io_mshrInfo_index ? _T_257_101_3 : _GEN_407;
  wire  _GEN_413 = 8'h66 == mshr_io_mshrInfo_index ? _T_257_102_1 : _GEN_409;
  wire  _GEN_414 = 8'h66 == mshr_io_mshrInfo_index ? _T_257_102_2 : _GEN_410;
  wire  _GEN_415 = 8'h66 == mshr_io_mshrInfo_index ? _T_257_102_3 : _GEN_411;
  wire  _GEN_417 = 8'h67 == mshr_io_mshrInfo_index ? _T_257_103_1 : _GEN_413;
  wire  _GEN_418 = 8'h67 == mshr_io_mshrInfo_index ? _T_257_103_2 : _GEN_414;
  wire  _GEN_419 = 8'h67 == mshr_io_mshrInfo_index ? _T_257_103_3 : _GEN_415;
  wire  _GEN_421 = 8'h68 == mshr_io_mshrInfo_index ? _T_257_104_1 : _GEN_417;
  wire  _GEN_422 = 8'h68 == mshr_io_mshrInfo_index ? _T_257_104_2 : _GEN_418;
  wire  _GEN_423 = 8'h68 == mshr_io_mshrInfo_index ? _T_257_104_3 : _GEN_419;
  wire  _GEN_425 = 8'h69 == mshr_io_mshrInfo_index ? _T_257_105_1 : _GEN_421;
  wire  _GEN_426 = 8'h69 == mshr_io_mshrInfo_index ? _T_257_105_2 : _GEN_422;
  wire  _GEN_427 = 8'h69 == mshr_io_mshrInfo_index ? _T_257_105_3 : _GEN_423;
  wire  _GEN_429 = 8'h6a == mshr_io_mshrInfo_index ? _T_257_106_1 : _GEN_425;
  wire  _GEN_430 = 8'h6a == mshr_io_mshrInfo_index ? _T_257_106_2 : _GEN_426;
  wire  _GEN_431 = 8'h6a == mshr_io_mshrInfo_index ? _T_257_106_3 : _GEN_427;
  wire  _GEN_433 = 8'h6b == mshr_io_mshrInfo_index ? _T_257_107_1 : _GEN_429;
  wire  _GEN_434 = 8'h6b == mshr_io_mshrInfo_index ? _T_257_107_2 : _GEN_430;
  wire  _GEN_435 = 8'h6b == mshr_io_mshrInfo_index ? _T_257_107_3 : _GEN_431;
  wire  _GEN_437 = 8'h6c == mshr_io_mshrInfo_index ? _T_257_108_1 : _GEN_433;
  wire  _GEN_438 = 8'h6c == mshr_io_mshrInfo_index ? _T_257_108_2 : _GEN_434;
  wire  _GEN_439 = 8'h6c == mshr_io_mshrInfo_index ? _T_257_108_3 : _GEN_435;
  wire  _GEN_441 = 8'h6d == mshr_io_mshrInfo_index ? _T_257_109_1 : _GEN_437;
  wire  _GEN_442 = 8'h6d == mshr_io_mshrInfo_index ? _T_257_109_2 : _GEN_438;
  wire  _GEN_443 = 8'h6d == mshr_io_mshrInfo_index ? _T_257_109_3 : _GEN_439;
  wire  _GEN_445 = 8'h6e == mshr_io_mshrInfo_index ? _T_257_110_1 : _GEN_441;
  wire  _GEN_446 = 8'h6e == mshr_io_mshrInfo_index ? _T_257_110_2 : _GEN_442;
  wire  _GEN_447 = 8'h6e == mshr_io_mshrInfo_index ? _T_257_110_3 : _GEN_443;
  wire  _GEN_449 = 8'h6f == mshr_io_mshrInfo_index ? _T_257_111_1 : _GEN_445;
  wire  _GEN_450 = 8'h6f == mshr_io_mshrInfo_index ? _T_257_111_2 : _GEN_446;
  wire  _GEN_451 = 8'h6f == mshr_io_mshrInfo_index ? _T_257_111_3 : _GEN_447;
  wire  _GEN_453 = 8'h70 == mshr_io_mshrInfo_index ? _T_257_112_1 : _GEN_449;
  wire  _GEN_454 = 8'h70 == mshr_io_mshrInfo_index ? _T_257_112_2 : _GEN_450;
  wire  _GEN_455 = 8'h70 == mshr_io_mshrInfo_index ? _T_257_112_3 : _GEN_451;
  wire  _GEN_457 = 8'h71 == mshr_io_mshrInfo_index ? _T_257_113_1 : _GEN_453;
  wire  _GEN_458 = 8'h71 == mshr_io_mshrInfo_index ? _T_257_113_2 : _GEN_454;
  wire  _GEN_459 = 8'h71 == mshr_io_mshrInfo_index ? _T_257_113_3 : _GEN_455;
  wire  _GEN_461 = 8'h72 == mshr_io_mshrInfo_index ? _T_257_114_1 : _GEN_457;
  wire  _GEN_462 = 8'h72 == mshr_io_mshrInfo_index ? _T_257_114_2 : _GEN_458;
  wire  _GEN_463 = 8'h72 == mshr_io_mshrInfo_index ? _T_257_114_3 : _GEN_459;
  wire  _GEN_465 = 8'h73 == mshr_io_mshrInfo_index ? _T_257_115_1 : _GEN_461;
  wire  _GEN_466 = 8'h73 == mshr_io_mshrInfo_index ? _T_257_115_2 : _GEN_462;
  wire  _GEN_467 = 8'h73 == mshr_io_mshrInfo_index ? _T_257_115_3 : _GEN_463;
  wire  _GEN_469 = 8'h74 == mshr_io_mshrInfo_index ? _T_257_116_1 : _GEN_465;
  wire  _GEN_470 = 8'h74 == mshr_io_mshrInfo_index ? _T_257_116_2 : _GEN_466;
  wire  _GEN_471 = 8'h74 == mshr_io_mshrInfo_index ? _T_257_116_3 : _GEN_467;
  wire  _GEN_473 = 8'h75 == mshr_io_mshrInfo_index ? _T_257_117_1 : _GEN_469;
  wire  _GEN_474 = 8'h75 == mshr_io_mshrInfo_index ? _T_257_117_2 : _GEN_470;
  wire  _GEN_475 = 8'h75 == mshr_io_mshrInfo_index ? _T_257_117_3 : _GEN_471;
  wire  _GEN_477 = 8'h76 == mshr_io_mshrInfo_index ? _T_257_118_1 : _GEN_473;
  wire  _GEN_478 = 8'h76 == mshr_io_mshrInfo_index ? _T_257_118_2 : _GEN_474;
  wire  _GEN_479 = 8'h76 == mshr_io_mshrInfo_index ? _T_257_118_3 : _GEN_475;
  wire  _GEN_481 = 8'h77 == mshr_io_mshrInfo_index ? _T_257_119_1 : _GEN_477;
  wire  _GEN_482 = 8'h77 == mshr_io_mshrInfo_index ? _T_257_119_2 : _GEN_478;
  wire  _GEN_483 = 8'h77 == mshr_io_mshrInfo_index ? _T_257_119_3 : _GEN_479;
  wire  _GEN_485 = 8'h78 == mshr_io_mshrInfo_index ? _T_257_120_1 : _GEN_481;
  wire  _GEN_486 = 8'h78 == mshr_io_mshrInfo_index ? _T_257_120_2 : _GEN_482;
  wire  _GEN_487 = 8'h78 == mshr_io_mshrInfo_index ? _T_257_120_3 : _GEN_483;
  wire  _GEN_489 = 8'h79 == mshr_io_mshrInfo_index ? _T_257_121_1 : _GEN_485;
  wire  _GEN_490 = 8'h79 == mshr_io_mshrInfo_index ? _T_257_121_2 : _GEN_486;
  wire  _GEN_491 = 8'h79 == mshr_io_mshrInfo_index ? _T_257_121_3 : _GEN_487;
  wire  _GEN_493 = 8'h7a == mshr_io_mshrInfo_index ? _T_257_122_1 : _GEN_489;
  wire  _GEN_494 = 8'h7a == mshr_io_mshrInfo_index ? _T_257_122_2 : _GEN_490;
  wire  _GEN_495 = 8'h7a == mshr_io_mshrInfo_index ? _T_257_122_3 : _GEN_491;
  wire  _GEN_497 = 8'h7b == mshr_io_mshrInfo_index ? _T_257_123_1 : _GEN_493;
  wire  _GEN_498 = 8'h7b == mshr_io_mshrInfo_index ? _T_257_123_2 : _GEN_494;
  wire  _GEN_499 = 8'h7b == mshr_io_mshrInfo_index ? _T_257_123_3 : _GEN_495;
  wire  _GEN_501 = 8'h7c == mshr_io_mshrInfo_index ? _T_257_124_1 : _GEN_497;
  wire  _GEN_502 = 8'h7c == mshr_io_mshrInfo_index ? _T_257_124_2 : _GEN_498;
  wire  _GEN_503 = 8'h7c == mshr_io_mshrInfo_index ? _T_257_124_3 : _GEN_499;
  wire  _GEN_505 = 8'h7d == mshr_io_mshrInfo_index ? _T_257_125_1 : _GEN_501;
  wire  _GEN_506 = 8'h7d == mshr_io_mshrInfo_index ? _T_257_125_2 : _GEN_502;
  wire  _GEN_507 = 8'h7d == mshr_io_mshrInfo_index ? _T_257_125_3 : _GEN_503;
  wire  _GEN_509 = 8'h7e == mshr_io_mshrInfo_index ? _T_257_126_1 : _GEN_505;
  wire  _GEN_510 = 8'h7e == mshr_io_mshrInfo_index ? _T_257_126_2 : _GEN_506;
  wire  _GEN_511 = 8'h7e == mshr_io_mshrInfo_index ? _T_257_126_3 : _GEN_507;
  wire  _GEN_513 = 8'h7f == mshr_io_mshrInfo_index ? _T_257_127_1 : _GEN_509;
  wire  _GEN_514 = 8'h7f == mshr_io_mshrInfo_index ? _T_257_127_2 : _GEN_510;
  wire  _GEN_515 = 8'h7f == mshr_io_mshrInfo_index ? _T_257_127_3 : _GEN_511;
  wire  _GEN_517 = 8'h80 == mshr_io_mshrInfo_index ? _T_257_128_1 : _GEN_513;
  wire  _GEN_518 = 8'h80 == mshr_io_mshrInfo_index ? _T_257_128_2 : _GEN_514;
  wire  _GEN_519 = 8'h80 == mshr_io_mshrInfo_index ? _T_257_128_3 : _GEN_515;
  wire  _GEN_521 = 8'h81 == mshr_io_mshrInfo_index ? _T_257_129_1 : _GEN_517;
  wire  _GEN_522 = 8'h81 == mshr_io_mshrInfo_index ? _T_257_129_2 : _GEN_518;
  wire  _GEN_523 = 8'h81 == mshr_io_mshrInfo_index ? _T_257_129_3 : _GEN_519;
  wire  _GEN_525 = 8'h82 == mshr_io_mshrInfo_index ? _T_257_130_1 : _GEN_521;
  wire  _GEN_526 = 8'h82 == mshr_io_mshrInfo_index ? _T_257_130_2 : _GEN_522;
  wire  _GEN_527 = 8'h82 == mshr_io_mshrInfo_index ? _T_257_130_3 : _GEN_523;
  wire  _GEN_529 = 8'h83 == mshr_io_mshrInfo_index ? _T_257_131_1 : _GEN_525;
  wire  _GEN_530 = 8'h83 == mshr_io_mshrInfo_index ? _T_257_131_2 : _GEN_526;
  wire  _GEN_531 = 8'h83 == mshr_io_mshrInfo_index ? _T_257_131_3 : _GEN_527;
  wire  _GEN_533 = 8'h84 == mshr_io_mshrInfo_index ? _T_257_132_1 : _GEN_529;
  wire  _GEN_534 = 8'h84 == mshr_io_mshrInfo_index ? _T_257_132_2 : _GEN_530;
  wire  _GEN_535 = 8'h84 == mshr_io_mshrInfo_index ? _T_257_132_3 : _GEN_531;
  wire  _GEN_537 = 8'h85 == mshr_io_mshrInfo_index ? _T_257_133_1 : _GEN_533;
  wire  _GEN_538 = 8'h85 == mshr_io_mshrInfo_index ? _T_257_133_2 : _GEN_534;
  wire  _GEN_539 = 8'h85 == mshr_io_mshrInfo_index ? _T_257_133_3 : _GEN_535;
  wire  _GEN_541 = 8'h86 == mshr_io_mshrInfo_index ? _T_257_134_1 : _GEN_537;
  wire  _GEN_542 = 8'h86 == mshr_io_mshrInfo_index ? _T_257_134_2 : _GEN_538;
  wire  _GEN_543 = 8'h86 == mshr_io_mshrInfo_index ? _T_257_134_3 : _GEN_539;
  wire  _GEN_545 = 8'h87 == mshr_io_mshrInfo_index ? _T_257_135_1 : _GEN_541;
  wire  _GEN_546 = 8'h87 == mshr_io_mshrInfo_index ? _T_257_135_2 : _GEN_542;
  wire  _GEN_547 = 8'h87 == mshr_io_mshrInfo_index ? _T_257_135_3 : _GEN_543;
  wire  _GEN_549 = 8'h88 == mshr_io_mshrInfo_index ? _T_257_136_1 : _GEN_545;
  wire  _GEN_550 = 8'h88 == mshr_io_mshrInfo_index ? _T_257_136_2 : _GEN_546;
  wire  _GEN_551 = 8'h88 == mshr_io_mshrInfo_index ? _T_257_136_3 : _GEN_547;
  wire  _GEN_553 = 8'h89 == mshr_io_mshrInfo_index ? _T_257_137_1 : _GEN_549;
  wire  _GEN_554 = 8'h89 == mshr_io_mshrInfo_index ? _T_257_137_2 : _GEN_550;
  wire  _GEN_555 = 8'h89 == mshr_io_mshrInfo_index ? _T_257_137_3 : _GEN_551;
  wire  _GEN_557 = 8'h8a == mshr_io_mshrInfo_index ? _T_257_138_1 : _GEN_553;
  wire  _GEN_558 = 8'h8a == mshr_io_mshrInfo_index ? _T_257_138_2 : _GEN_554;
  wire  _GEN_559 = 8'h8a == mshr_io_mshrInfo_index ? _T_257_138_3 : _GEN_555;
  wire  _GEN_561 = 8'h8b == mshr_io_mshrInfo_index ? _T_257_139_1 : _GEN_557;
  wire  _GEN_562 = 8'h8b == mshr_io_mshrInfo_index ? _T_257_139_2 : _GEN_558;
  wire  _GEN_563 = 8'h8b == mshr_io_mshrInfo_index ? _T_257_139_3 : _GEN_559;
  wire  _GEN_565 = 8'h8c == mshr_io_mshrInfo_index ? _T_257_140_1 : _GEN_561;
  wire  _GEN_566 = 8'h8c == mshr_io_mshrInfo_index ? _T_257_140_2 : _GEN_562;
  wire  _GEN_567 = 8'h8c == mshr_io_mshrInfo_index ? _T_257_140_3 : _GEN_563;
  wire  _GEN_569 = 8'h8d == mshr_io_mshrInfo_index ? _T_257_141_1 : _GEN_565;
  wire  _GEN_570 = 8'h8d == mshr_io_mshrInfo_index ? _T_257_141_2 : _GEN_566;
  wire  _GEN_571 = 8'h8d == mshr_io_mshrInfo_index ? _T_257_141_3 : _GEN_567;
  wire  _GEN_573 = 8'h8e == mshr_io_mshrInfo_index ? _T_257_142_1 : _GEN_569;
  wire  _GEN_574 = 8'h8e == mshr_io_mshrInfo_index ? _T_257_142_2 : _GEN_570;
  wire  _GEN_575 = 8'h8e == mshr_io_mshrInfo_index ? _T_257_142_3 : _GEN_571;
  wire  _GEN_577 = 8'h8f == mshr_io_mshrInfo_index ? _T_257_143_1 : _GEN_573;
  wire  _GEN_578 = 8'h8f == mshr_io_mshrInfo_index ? _T_257_143_2 : _GEN_574;
  wire  _GEN_579 = 8'h8f == mshr_io_mshrInfo_index ? _T_257_143_3 : _GEN_575;
  wire  _GEN_581 = 8'h90 == mshr_io_mshrInfo_index ? _T_257_144_1 : _GEN_577;
  wire  _GEN_582 = 8'h90 == mshr_io_mshrInfo_index ? _T_257_144_2 : _GEN_578;
  wire  _GEN_583 = 8'h90 == mshr_io_mshrInfo_index ? _T_257_144_3 : _GEN_579;
  wire  _GEN_585 = 8'h91 == mshr_io_mshrInfo_index ? _T_257_145_1 : _GEN_581;
  wire  _GEN_586 = 8'h91 == mshr_io_mshrInfo_index ? _T_257_145_2 : _GEN_582;
  wire  _GEN_587 = 8'h91 == mshr_io_mshrInfo_index ? _T_257_145_3 : _GEN_583;
  wire  _GEN_589 = 8'h92 == mshr_io_mshrInfo_index ? _T_257_146_1 : _GEN_585;
  wire  _GEN_590 = 8'h92 == mshr_io_mshrInfo_index ? _T_257_146_2 : _GEN_586;
  wire  _GEN_591 = 8'h92 == mshr_io_mshrInfo_index ? _T_257_146_3 : _GEN_587;
  wire  _GEN_593 = 8'h93 == mshr_io_mshrInfo_index ? _T_257_147_1 : _GEN_589;
  wire  _GEN_594 = 8'h93 == mshr_io_mshrInfo_index ? _T_257_147_2 : _GEN_590;
  wire  _GEN_595 = 8'h93 == mshr_io_mshrInfo_index ? _T_257_147_3 : _GEN_591;
  wire  _GEN_597 = 8'h94 == mshr_io_mshrInfo_index ? _T_257_148_1 : _GEN_593;
  wire  _GEN_598 = 8'h94 == mshr_io_mshrInfo_index ? _T_257_148_2 : _GEN_594;
  wire  _GEN_599 = 8'h94 == mshr_io_mshrInfo_index ? _T_257_148_3 : _GEN_595;
  wire  _GEN_601 = 8'h95 == mshr_io_mshrInfo_index ? _T_257_149_1 : _GEN_597;
  wire  _GEN_602 = 8'h95 == mshr_io_mshrInfo_index ? _T_257_149_2 : _GEN_598;
  wire  _GEN_603 = 8'h95 == mshr_io_mshrInfo_index ? _T_257_149_3 : _GEN_599;
  wire  _GEN_605 = 8'h96 == mshr_io_mshrInfo_index ? _T_257_150_1 : _GEN_601;
  wire  _GEN_606 = 8'h96 == mshr_io_mshrInfo_index ? _T_257_150_2 : _GEN_602;
  wire  _GEN_607 = 8'h96 == mshr_io_mshrInfo_index ? _T_257_150_3 : _GEN_603;
  wire  _GEN_609 = 8'h97 == mshr_io_mshrInfo_index ? _T_257_151_1 : _GEN_605;
  wire  _GEN_610 = 8'h97 == mshr_io_mshrInfo_index ? _T_257_151_2 : _GEN_606;
  wire  _GEN_611 = 8'h97 == mshr_io_mshrInfo_index ? _T_257_151_3 : _GEN_607;
  wire  _GEN_613 = 8'h98 == mshr_io_mshrInfo_index ? _T_257_152_1 : _GEN_609;
  wire  _GEN_614 = 8'h98 == mshr_io_mshrInfo_index ? _T_257_152_2 : _GEN_610;
  wire  _GEN_615 = 8'h98 == mshr_io_mshrInfo_index ? _T_257_152_3 : _GEN_611;
  wire  _GEN_617 = 8'h99 == mshr_io_mshrInfo_index ? _T_257_153_1 : _GEN_613;
  wire  _GEN_618 = 8'h99 == mshr_io_mshrInfo_index ? _T_257_153_2 : _GEN_614;
  wire  _GEN_619 = 8'h99 == mshr_io_mshrInfo_index ? _T_257_153_3 : _GEN_615;
  wire  _GEN_621 = 8'h9a == mshr_io_mshrInfo_index ? _T_257_154_1 : _GEN_617;
  wire  _GEN_622 = 8'h9a == mshr_io_mshrInfo_index ? _T_257_154_2 : _GEN_618;
  wire  _GEN_623 = 8'h9a == mshr_io_mshrInfo_index ? _T_257_154_3 : _GEN_619;
  wire  _GEN_625 = 8'h9b == mshr_io_mshrInfo_index ? _T_257_155_1 : _GEN_621;
  wire  _GEN_626 = 8'h9b == mshr_io_mshrInfo_index ? _T_257_155_2 : _GEN_622;
  wire  _GEN_627 = 8'h9b == mshr_io_mshrInfo_index ? _T_257_155_3 : _GEN_623;
  wire  _GEN_629 = 8'h9c == mshr_io_mshrInfo_index ? _T_257_156_1 : _GEN_625;
  wire  _GEN_630 = 8'h9c == mshr_io_mshrInfo_index ? _T_257_156_2 : _GEN_626;
  wire  _GEN_631 = 8'h9c == mshr_io_mshrInfo_index ? _T_257_156_3 : _GEN_627;
  wire  _GEN_633 = 8'h9d == mshr_io_mshrInfo_index ? _T_257_157_1 : _GEN_629;
  wire  _GEN_634 = 8'h9d == mshr_io_mshrInfo_index ? _T_257_157_2 : _GEN_630;
  wire  _GEN_635 = 8'h9d == mshr_io_mshrInfo_index ? _T_257_157_3 : _GEN_631;
  wire  _GEN_637 = 8'h9e == mshr_io_mshrInfo_index ? _T_257_158_1 : _GEN_633;
  wire  _GEN_638 = 8'h9e == mshr_io_mshrInfo_index ? _T_257_158_2 : _GEN_634;
  wire  _GEN_639 = 8'h9e == mshr_io_mshrInfo_index ? _T_257_158_3 : _GEN_635;
  wire  _GEN_641 = 8'h9f == mshr_io_mshrInfo_index ? _T_257_159_1 : _GEN_637;
  wire  _GEN_642 = 8'h9f == mshr_io_mshrInfo_index ? _T_257_159_2 : _GEN_638;
  wire  _GEN_643 = 8'h9f == mshr_io_mshrInfo_index ? _T_257_159_3 : _GEN_639;
  wire  _GEN_645 = 8'ha0 == mshr_io_mshrInfo_index ? _T_257_160_1 : _GEN_641;
  wire  _GEN_646 = 8'ha0 == mshr_io_mshrInfo_index ? _T_257_160_2 : _GEN_642;
  wire  _GEN_647 = 8'ha0 == mshr_io_mshrInfo_index ? _T_257_160_3 : _GEN_643;
  wire  _GEN_649 = 8'ha1 == mshr_io_mshrInfo_index ? _T_257_161_1 : _GEN_645;
  wire  _GEN_650 = 8'ha1 == mshr_io_mshrInfo_index ? _T_257_161_2 : _GEN_646;
  wire  _GEN_651 = 8'ha1 == mshr_io_mshrInfo_index ? _T_257_161_3 : _GEN_647;
  wire  _GEN_653 = 8'ha2 == mshr_io_mshrInfo_index ? _T_257_162_1 : _GEN_649;
  wire  _GEN_654 = 8'ha2 == mshr_io_mshrInfo_index ? _T_257_162_2 : _GEN_650;
  wire  _GEN_655 = 8'ha2 == mshr_io_mshrInfo_index ? _T_257_162_3 : _GEN_651;
  wire  _GEN_657 = 8'ha3 == mshr_io_mshrInfo_index ? _T_257_163_1 : _GEN_653;
  wire  _GEN_658 = 8'ha3 == mshr_io_mshrInfo_index ? _T_257_163_2 : _GEN_654;
  wire  _GEN_659 = 8'ha3 == mshr_io_mshrInfo_index ? _T_257_163_3 : _GEN_655;
  wire  _GEN_661 = 8'ha4 == mshr_io_mshrInfo_index ? _T_257_164_1 : _GEN_657;
  wire  _GEN_662 = 8'ha4 == mshr_io_mshrInfo_index ? _T_257_164_2 : _GEN_658;
  wire  _GEN_663 = 8'ha4 == mshr_io_mshrInfo_index ? _T_257_164_3 : _GEN_659;
  wire  _GEN_665 = 8'ha5 == mshr_io_mshrInfo_index ? _T_257_165_1 : _GEN_661;
  wire  _GEN_666 = 8'ha5 == mshr_io_mshrInfo_index ? _T_257_165_2 : _GEN_662;
  wire  _GEN_667 = 8'ha5 == mshr_io_mshrInfo_index ? _T_257_165_3 : _GEN_663;
  wire  _GEN_669 = 8'ha6 == mshr_io_mshrInfo_index ? _T_257_166_1 : _GEN_665;
  wire  _GEN_670 = 8'ha6 == mshr_io_mshrInfo_index ? _T_257_166_2 : _GEN_666;
  wire  _GEN_671 = 8'ha6 == mshr_io_mshrInfo_index ? _T_257_166_3 : _GEN_667;
  wire  _GEN_673 = 8'ha7 == mshr_io_mshrInfo_index ? _T_257_167_1 : _GEN_669;
  wire  _GEN_674 = 8'ha7 == mshr_io_mshrInfo_index ? _T_257_167_2 : _GEN_670;
  wire  _GEN_675 = 8'ha7 == mshr_io_mshrInfo_index ? _T_257_167_3 : _GEN_671;
  wire  _GEN_677 = 8'ha8 == mshr_io_mshrInfo_index ? _T_257_168_1 : _GEN_673;
  wire  _GEN_678 = 8'ha8 == mshr_io_mshrInfo_index ? _T_257_168_2 : _GEN_674;
  wire  _GEN_679 = 8'ha8 == mshr_io_mshrInfo_index ? _T_257_168_3 : _GEN_675;
  wire  _GEN_681 = 8'ha9 == mshr_io_mshrInfo_index ? _T_257_169_1 : _GEN_677;
  wire  _GEN_682 = 8'ha9 == mshr_io_mshrInfo_index ? _T_257_169_2 : _GEN_678;
  wire  _GEN_683 = 8'ha9 == mshr_io_mshrInfo_index ? _T_257_169_3 : _GEN_679;
  wire  _GEN_685 = 8'haa == mshr_io_mshrInfo_index ? _T_257_170_1 : _GEN_681;
  wire  _GEN_686 = 8'haa == mshr_io_mshrInfo_index ? _T_257_170_2 : _GEN_682;
  wire  _GEN_687 = 8'haa == mshr_io_mshrInfo_index ? _T_257_170_3 : _GEN_683;
  wire  _GEN_689 = 8'hab == mshr_io_mshrInfo_index ? _T_257_171_1 : _GEN_685;
  wire  _GEN_690 = 8'hab == mshr_io_mshrInfo_index ? _T_257_171_2 : _GEN_686;
  wire  _GEN_691 = 8'hab == mshr_io_mshrInfo_index ? _T_257_171_3 : _GEN_687;
  wire  _GEN_693 = 8'hac == mshr_io_mshrInfo_index ? _T_257_172_1 : _GEN_689;
  wire  _GEN_694 = 8'hac == mshr_io_mshrInfo_index ? _T_257_172_2 : _GEN_690;
  wire  _GEN_695 = 8'hac == mshr_io_mshrInfo_index ? _T_257_172_3 : _GEN_691;
  wire  _GEN_697 = 8'had == mshr_io_mshrInfo_index ? _T_257_173_1 : _GEN_693;
  wire  _GEN_698 = 8'had == mshr_io_mshrInfo_index ? _T_257_173_2 : _GEN_694;
  wire  _GEN_699 = 8'had == mshr_io_mshrInfo_index ? _T_257_173_3 : _GEN_695;
  wire  _GEN_701 = 8'hae == mshr_io_mshrInfo_index ? _T_257_174_1 : _GEN_697;
  wire  _GEN_702 = 8'hae == mshr_io_mshrInfo_index ? _T_257_174_2 : _GEN_698;
  wire  _GEN_703 = 8'hae == mshr_io_mshrInfo_index ? _T_257_174_3 : _GEN_699;
  wire  _GEN_705 = 8'haf == mshr_io_mshrInfo_index ? _T_257_175_1 : _GEN_701;
  wire  _GEN_706 = 8'haf == mshr_io_mshrInfo_index ? _T_257_175_2 : _GEN_702;
  wire  _GEN_707 = 8'haf == mshr_io_mshrInfo_index ? _T_257_175_3 : _GEN_703;
  wire  _GEN_709 = 8'hb0 == mshr_io_mshrInfo_index ? _T_257_176_1 : _GEN_705;
  wire  _GEN_710 = 8'hb0 == mshr_io_mshrInfo_index ? _T_257_176_2 : _GEN_706;
  wire  _GEN_711 = 8'hb0 == mshr_io_mshrInfo_index ? _T_257_176_3 : _GEN_707;
  wire  _GEN_713 = 8'hb1 == mshr_io_mshrInfo_index ? _T_257_177_1 : _GEN_709;
  wire  _GEN_714 = 8'hb1 == mshr_io_mshrInfo_index ? _T_257_177_2 : _GEN_710;
  wire  _GEN_715 = 8'hb1 == mshr_io_mshrInfo_index ? _T_257_177_3 : _GEN_711;
  wire  _GEN_717 = 8'hb2 == mshr_io_mshrInfo_index ? _T_257_178_1 : _GEN_713;
  wire  _GEN_718 = 8'hb2 == mshr_io_mshrInfo_index ? _T_257_178_2 : _GEN_714;
  wire  _GEN_719 = 8'hb2 == mshr_io_mshrInfo_index ? _T_257_178_3 : _GEN_715;
  wire  _GEN_721 = 8'hb3 == mshr_io_mshrInfo_index ? _T_257_179_1 : _GEN_717;
  wire  _GEN_722 = 8'hb3 == mshr_io_mshrInfo_index ? _T_257_179_2 : _GEN_718;
  wire  _GEN_723 = 8'hb3 == mshr_io_mshrInfo_index ? _T_257_179_3 : _GEN_719;
  wire  _GEN_725 = 8'hb4 == mshr_io_mshrInfo_index ? _T_257_180_1 : _GEN_721;
  wire  _GEN_726 = 8'hb4 == mshr_io_mshrInfo_index ? _T_257_180_2 : _GEN_722;
  wire  _GEN_727 = 8'hb4 == mshr_io_mshrInfo_index ? _T_257_180_3 : _GEN_723;
  wire  _GEN_729 = 8'hb5 == mshr_io_mshrInfo_index ? _T_257_181_1 : _GEN_725;
  wire  _GEN_730 = 8'hb5 == mshr_io_mshrInfo_index ? _T_257_181_2 : _GEN_726;
  wire  _GEN_731 = 8'hb5 == mshr_io_mshrInfo_index ? _T_257_181_3 : _GEN_727;
  wire  _GEN_733 = 8'hb6 == mshr_io_mshrInfo_index ? _T_257_182_1 : _GEN_729;
  wire  _GEN_734 = 8'hb6 == mshr_io_mshrInfo_index ? _T_257_182_2 : _GEN_730;
  wire  _GEN_735 = 8'hb6 == mshr_io_mshrInfo_index ? _T_257_182_3 : _GEN_731;
  wire  _GEN_737 = 8'hb7 == mshr_io_mshrInfo_index ? _T_257_183_1 : _GEN_733;
  wire  _GEN_738 = 8'hb7 == mshr_io_mshrInfo_index ? _T_257_183_2 : _GEN_734;
  wire  _GEN_739 = 8'hb7 == mshr_io_mshrInfo_index ? _T_257_183_3 : _GEN_735;
  wire  _GEN_741 = 8'hb8 == mshr_io_mshrInfo_index ? _T_257_184_1 : _GEN_737;
  wire  _GEN_742 = 8'hb8 == mshr_io_mshrInfo_index ? _T_257_184_2 : _GEN_738;
  wire  _GEN_743 = 8'hb8 == mshr_io_mshrInfo_index ? _T_257_184_3 : _GEN_739;
  wire  _GEN_745 = 8'hb9 == mshr_io_mshrInfo_index ? _T_257_185_1 : _GEN_741;
  wire  _GEN_746 = 8'hb9 == mshr_io_mshrInfo_index ? _T_257_185_2 : _GEN_742;
  wire  _GEN_747 = 8'hb9 == mshr_io_mshrInfo_index ? _T_257_185_3 : _GEN_743;
  wire  _GEN_749 = 8'hba == mshr_io_mshrInfo_index ? _T_257_186_1 : _GEN_745;
  wire  _GEN_750 = 8'hba == mshr_io_mshrInfo_index ? _T_257_186_2 : _GEN_746;
  wire  _GEN_751 = 8'hba == mshr_io_mshrInfo_index ? _T_257_186_3 : _GEN_747;
  wire  _GEN_753 = 8'hbb == mshr_io_mshrInfo_index ? _T_257_187_1 : _GEN_749;
  wire  _GEN_754 = 8'hbb == mshr_io_mshrInfo_index ? _T_257_187_2 : _GEN_750;
  wire  _GEN_755 = 8'hbb == mshr_io_mshrInfo_index ? _T_257_187_3 : _GEN_751;
  wire  _GEN_757 = 8'hbc == mshr_io_mshrInfo_index ? _T_257_188_1 : _GEN_753;
  wire  _GEN_758 = 8'hbc == mshr_io_mshrInfo_index ? _T_257_188_2 : _GEN_754;
  wire  _GEN_759 = 8'hbc == mshr_io_mshrInfo_index ? _T_257_188_3 : _GEN_755;
  wire  _GEN_761 = 8'hbd == mshr_io_mshrInfo_index ? _T_257_189_1 : _GEN_757;
  wire  _GEN_762 = 8'hbd == mshr_io_mshrInfo_index ? _T_257_189_2 : _GEN_758;
  wire  _GEN_763 = 8'hbd == mshr_io_mshrInfo_index ? _T_257_189_3 : _GEN_759;
  wire  _GEN_765 = 8'hbe == mshr_io_mshrInfo_index ? _T_257_190_1 : _GEN_761;
  wire  _GEN_766 = 8'hbe == mshr_io_mshrInfo_index ? _T_257_190_2 : _GEN_762;
  wire  _GEN_767 = 8'hbe == mshr_io_mshrInfo_index ? _T_257_190_3 : _GEN_763;
  wire  _GEN_769 = 8'hbf == mshr_io_mshrInfo_index ? _T_257_191_1 : _GEN_765;
  wire  _GEN_770 = 8'hbf == mshr_io_mshrInfo_index ? _T_257_191_2 : _GEN_766;
  wire  _GEN_771 = 8'hbf == mshr_io_mshrInfo_index ? _T_257_191_3 : _GEN_767;
  wire  _GEN_773 = 8'hc0 == mshr_io_mshrInfo_index ? _T_257_192_1 : _GEN_769;
  wire  _GEN_774 = 8'hc0 == mshr_io_mshrInfo_index ? _T_257_192_2 : _GEN_770;
  wire  _GEN_775 = 8'hc0 == mshr_io_mshrInfo_index ? _T_257_192_3 : _GEN_771;
  wire  _GEN_777 = 8'hc1 == mshr_io_mshrInfo_index ? _T_257_193_1 : _GEN_773;
  wire  _GEN_778 = 8'hc1 == mshr_io_mshrInfo_index ? _T_257_193_2 : _GEN_774;
  wire  _GEN_779 = 8'hc1 == mshr_io_mshrInfo_index ? _T_257_193_3 : _GEN_775;
  wire  _GEN_781 = 8'hc2 == mshr_io_mshrInfo_index ? _T_257_194_1 : _GEN_777;
  wire  _GEN_782 = 8'hc2 == mshr_io_mshrInfo_index ? _T_257_194_2 : _GEN_778;
  wire  _GEN_783 = 8'hc2 == mshr_io_mshrInfo_index ? _T_257_194_3 : _GEN_779;
  wire  _GEN_785 = 8'hc3 == mshr_io_mshrInfo_index ? _T_257_195_1 : _GEN_781;
  wire  _GEN_786 = 8'hc3 == mshr_io_mshrInfo_index ? _T_257_195_2 : _GEN_782;
  wire  _GEN_787 = 8'hc3 == mshr_io_mshrInfo_index ? _T_257_195_3 : _GEN_783;
  wire  _GEN_789 = 8'hc4 == mshr_io_mshrInfo_index ? _T_257_196_1 : _GEN_785;
  wire  _GEN_790 = 8'hc4 == mshr_io_mshrInfo_index ? _T_257_196_2 : _GEN_786;
  wire  _GEN_791 = 8'hc4 == mshr_io_mshrInfo_index ? _T_257_196_3 : _GEN_787;
  wire  _GEN_793 = 8'hc5 == mshr_io_mshrInfo_index ? _T_257_197_1 : _GEN_789;
  wire  _GEN_794 = 8'hc5 == mshr_io_mshrInfo_index ? _T_257_197_2 : _GEN_790;
  wire  _GEN_795 = 8'hc5 == mshr_io_mshrInfo_index ? _T_257_197_3 : _GEN_791;
  wire  _GEN_797 = 8'hc6 == mshr_io_mshrInfo_index ? _T_257_198_1 : _GEN_793;
  wire  _GEN_798 = 8'hc6 == mshr_io_mshrInfo_index ? _T_257_198_2 : _GEN_794;
  wire  _GEN_799 = 8'hc6 == mshr_io_mshrInfo_index ? _T_257_198_3 : _GEN_795;
  wire  _GEN_801 = 8'hc7 == mshr_io_mshrInfo_index ? _T_257_199_1 : _GEN_797;
  wire  _GEN_802 = 8'hc7 == mshr_io_mshrInfo_index ? _T_257_199_2 : _GEN_798;
  wire  _GEN_803 = 8'hc7 == mshr_io_mshrInfo_index ? _T_257_199_3 : _GEN_799;
  wire  _GEN_805 = 8'hc8 == mshr_io_mshrInfo_index ? _T_257_200_1 : _GEN_801;
  wire  _GEN_806 = 8'hc8 == mshr_io_mshrInfo_index ? _T_257_200_2 : _GEN_802;
  wire  _GEN_807 = 8'hc8 == mshr_io_mshrInfo_index ? _T_257_200_3 : _GEN_803;
  wire  _GEN_809 = 8'hc9 == mshr_io_mshrInfo_index ? _T_257_201_1 : _GEN_805;
  wire  _GEN_810 = 8'hc9 == mshr_io_mshrInfo_index ? _T_257_201_2 : _GEN_806;
  wire  _GEN_811 = 8'hc9 == mshr_io_mshrInfo_index ? _T_257_201_3 : _GEN_807;
  wire  _GEN_813 = 8'hca == mshr_io_mshrInfo_index ? _T_257_202_1 : _GEN_809;
  wire  _GEN_814 = 8'hca == mshr_io_mshrInfo_index ? _T_257_202_2 : _GEN_810;
  wire  _GEN_815 = 8'hca == mshr_io_mshrInfo_index ? _T_257_202_3 : _GEN_811;
  wire  _GEN_817 = 8'hcb == mshr_io_mshrInfo_index ? _T_257_203_1 : _GEN_813;
  wire  _GEN_818 = 8'hcb == mshr_io_mshrInfo_index ? _T_257_203_2 : _GEN_814;
  wire  _GEN_819 = 8'hcb == mshr_io_mshrInfo_index ? _T_257_203_3 : _GEN_815;
  wire  _GEN_821 = 8'hcc == mshr_io_mshrInfo_index ? _T_257_204_1 : _GEN_817;
  wire  _GEN_822 = 8'hcc == mshr_io_mshrInfo_index ? _T_257_204_2 : _GEN_818;
  wire  _GEN_823 = 8'hcc == mshr_io_mshrInfo_index ? _T_257_204_3 : _GEN_819;
  wire  _GEN_825 = 8'hcd == mshr_io_mshrInfo_index ? _T_257_205_1 : _GEN_821;
  wire  _GEN_826 = 8'hcd == mshr_io_mshrInfo_index ? _T_257_205_2 : _GEN_822;
  wire  _GEN_827 = 8'hcd == mshr_io_mshrInfo_index ? _T_257_205_3 : _GEN_823;
  wire  _GEN_829 = 8'hce == mshr_io_mshrInfo_index ? _T_257_206_1 : _GEN_825;
  wire  _GEN_830 = 8'hce == mshr_io_mshrInfo_index ? _T_257_206_2 : _GEN_826;
  wire  _GEN_831 = 8'hce == mshr_io_mshrInfo_index ? _T_257_206_3 : _GEN_827;
  wire  _GEN_833 = 8'hcf == mshr_io_mshrInfo_index ? _T_257_207_1 : _GEN_829;
  wire  _GEN_834 = 8'hcf == mshr_io_mshrInfo_index ? _T_257_207_2 : _GEN_830;
  wire  _GEN_835 = 8'hcf == mshr_io_mshrInfo_index ? _T_257_207_3 : _GEN_831;
  wire  _GEN_837 = 8'hd0 == mshr_io_mshrInfo_index ? _T_257_208_1 : _GEN_833;
  wire  _GEN_838 = 8'hd0 == mshr_io_mshrInfo_index ? _T_257_208_2 : _GEN_834;
  wire  _GEN_839 = 8'hd0 == mshr_io_mshrInfo_index ? _T_257_208_3 : _GEN_835;
  wire  _GEN_841 = 8'hd1 == mshr_io_mshrInfo_index ? _T_257_209_1 : _GEN_837;
  wire  _GEN_842 = 8'hd1 == mshr_io_mshrInfo_index ? _T_257_209_2 : _GEN_838;
  wire  _GEN_843 = 8'hd1 == mshr_io_mshrInfo_index ? _T_257_209_3 : _GEN_839;
  wire  _GEN_845 = 8'hd2 == mshr_io_mshrInfo_index ? _T_257_210_1 : _GEN_841;
  wire  _GEN_846 = 8'hd2 == mshr_io_mshrInfo_index ? _T_257_210_2 : _GEN_842;
  wire  _GEN_847 = 8'hd2 == mshr_io_mshrInfo_index ? _T_257_210_3 : _GEN_843;
  wire  _GEN_849 = 8'hd3 == mshr_io_mshrInfo_index ? _T_257_211_1 : _GEN_845;
  wire  _GEN_850 = 8'hd3 == mshr_io_mshrInfo_index ? _T_257_211_2 : _GEN_846;
  wire  _GEN_851 = 8'hd3 == mshr_io_mshrInfo_index ? _T_257_211_3 : _GEN_847;
  wire  _GEN_853 = 8'hd4 == mshr_io_mshrInfo_index ? _T_257_212_1 : _GEN_849;
  wire  _GEN_854 = 8'hd4 == mshr_io_mshrInfo_index ? _T_257_212_2 : _GEN_850;
  wire  _GEN_855 = 8'hd4 == mshr_io_mshrInfo_index ? _T_257_212_3 : _GEN_851;
  wire  _GEN_857 = 8'hd5 == mshr_io_mshrInfo_index ? _T_257_213_1 : _GEN_853;
  wire  _GEN_858 = 8'hd5 == mshr_io_mshrInfo_index ? _T_257_213_2 : _GEN_854;
  wire  _GEN_859 = 8'hd5 == mshr_io_mshrInfo_index ? _T_257_213_3 : _GEN_855;
  wire  _GEN_861 = 8'hd6 == mshr_io_mshrInfo_index ? _T_257_214_1 : _GEN_857;
  wire  _GEN_862 = 8'hd6 == mshr_io_mshrInfo_index ? _T_257_214_2 : _GEN_858;
  wire  _GEN_863 = 8'hd6 == mshr_io_mshrInfo_index ? _T_257_214_3 : _GEN_859;
  wire  _GEN_865 = 8'hd7 == mshr_io_mshrInfo_index ? _T_257_215_1 : _GEN_861;
  wire  _GEN_866 = 8'hd7 == mshr_io_mshrInfo_index ? _T_257_215_2 : _GEN_862;
  wire  _GEN_867 = 8'hd7 == mshr_io_mshrInfo_index ? _T_257_215_3 : _GEN_863;
  wire  _GEN_869 = 8'hd8 == mshr_io_mshrInfo_index ? _T_257_216_1 : _GEN_865;
  wire  _GEN_870 = 8'hd8 == mshr_io_mshrInfo_index ? _T_257_216_2 : _GEN_866;
  wire  _GEN_871 = 8'hd8 == mshr_io_mshrInfo_index ? _T_257_216_3 : _GEN_867;
  wire  _GEN_873 = 8'hd9 == mshr_io_mshrInfo_index ? _T_257_217_1 : _GEN_869;
  wire  _GEN_874 = 8'hd9 == mshr_io_mshrInfo_index ? _T_257_217_2 : _GEN_870;
  wire  _GEN_875 = 8'hd9 == mshr_io_mshrInfo_index ? _T_257_217_3 : _GEN_871;
  wire  _GEN_877 = 8'hda == mshr_io_mshrInfo_index ? _T_257_218_1 : _GEN_873;
  wire  _GEN_878 = 8'hda == mshr_io_mshrInfo_index ? _T_257_218_2 : _GEN_874;
  wire  _GEN_879 = 8'hda == mshr_io_mshrInfo_index ? _T_257_218_3 : _GEN_875;
  wire  _GEN_881 = 8'hdb == mshr_io_mshrInfo_index ? _T_257_219_1 : _GEN_877;
  wire  _GEN_882 = 8'hdb == mshr_io_mshrInfo_index ? _T_257_219_2 : _GEN_878;
  wire  _GEN_883 = 8'hdb == mshr_io_mshrInfo_index ? _T_257_219_3 : _GEN_879;
  wire  _GEN_885 = 8'hdc == mshr_io_mshrInfo_index ? _T_257_220_1 : _GEN_881;
  wire  _GEN_886 = 8'hdc == mshr_io_mshrInfo_index ? _T_257_220_2 : _GEN_882;
  wire  _GEN_887 = 8'hdc == mshr_io_mshrInfo_index ? _T_257_220_3 : _GEN_883;
  wire  _GEN_889 = 8'hdd == mshr_io_mshrInfo_index ? _T_257_221_1 : _GEN_885;
  wire  _GEN_890 = 8'hdd == mshr_io_mshrInfo_index ? _T_257_221_2 : _GEN_886;
  wire  _GEN_891 = 8'hdd == mshr_io_mshrInfo_index ? _T_257_221_3 : _GEN_887;
  wire  _GEN_893 = 8'hde == mshr_io_mshrInfo_index ? _T_257_222_1 : _GEN_889;
  wire  _GEN_894 = 8'hde == mshr_io_mshrInfo_index ? _T_257_222_2 : _GEN_890;
  wire  _GEN_895 = 8'hde == mshr_io_mshrInfo_index ? _T_257_222_3 : _GEN_891;
  wire  _GEN_897 = 8'hdf == mshr_io_mshrInfo_index ? _T_257_223_1 : _GEN_893;
  wire  _GEN_898 = 8'hdf == mshr_io_mshrInfo_index ? _T_257_223_2 : _GEN_894;
  wire  _GEN_899 = 8'hdf == mshr_io_mshrInfo_index ? _T_257_223_3 : _GEN_895;
  wire  _GEN_901 = 8'he0 == mshr_io_mshrInfo_index ? _T_257_224_1 : _GEN_897;
  wire  _GEN_902 = 8'he0 == mshr_io_mshrInfo_index ? _T_257_224_2 : _GEN_898;
  wire  _GEN_903 = 8'he0 == mshr_io_mshrInfo_index ? _T_257_224_3 : _GEN_899;
  wire  _GEN_905 = 8'he1 == mshr_io_mshrInfo_index ? _T_257_225_1 : _GEN_901;
  wire  _GEN_906 = 8'he1 == mshr_io_mshrInfo_index ? _T_257_225_2 : _GEN_902;
  wire  _GEN_907 = 8'he1 == mshr_io_mshrInfo_index ? _T_257_225_3 : _GEN_903;
  wire  _GEN_909 = 8'he2 == mshr_io_mshrInfo_index ? _T_257_226_1 : _GEN_905;
  wire  _GEN_910 = 8'he2 == mshr_io_mshrInfo_index ? _T_257_226_2 : _GEN_906;
  wire  _GEN_911 = 8'he2 == mshr_io_mshrInfo_index ? _T_257_226_3 : _GEN_907;
  wire  _GEN_913 = 8'he3 == mshr_io_mshrInfo_index ? _T_257_227_1 : _GEN_909;
  wire  _GEN_914 = 8'he3 == mshr_io_mshrInfo_index ? _T_257_227_2 : _GEN_910;
  wire  _GEN_915 = 8'he3 == mshr_io_mshrInfo_index ? _T_257_227_3 : _GEN_911;
  wire  _GEN_917 = 8'he4 == mshr_io_mshrInfo_index ? _T_257_228_1 : _GEN_913;
  wire  _GEN_918 = 8'he4 == mshr_io_mshrInfo_index ? _T_257_228_2 : _GEN_914;
  wire  _GEN_919 = 8'he4 == mshr_io_mshrInfo_index ? _T_257_228_3 : _GEN_915;
  wire  _GEN_921 = 8'he5 == mshr_io_mshrInfo_index ? _T_257_229_1 : _GEN_917;
  wire  _GEN_922 = 8'he5 == mshr_io_mshrInfo_index ? _T_257_229_2 : _GEN_918;
  wire  _GEN_923 = 8'he5 == mshr_io_mshrInfo_index ? _T_257_229_3 : _GEN_919;
  wire  _GEN_925 = 8'he6 == mshr_io_mshrInfo_index ? _T_257_230_1 : _GEN_921;
  wire  _GEN_926 = 8'he6 == mshr_io_mshrInfo_index ? _T_257_230_2 : _GEN_922;
  wire  _GEN_927 = 8'he6 == mshr_io_mshrInfo_index ? _T_257_230_3 : _GEN_923;
  wire  _GEN_929 = 8'he7 == mshr_io_mshrInfo_index ? _T_257_231_1 : _GEN_925;
  wire  _GEN_930 = 8'he7 == mshr_io_mshrInfo_index ? _T_257_231_2 : _GEN_926;
  wire  _GEN_931 = 8'he7 == mshr_io_mshrInfo_index ? _T_257_231_3 : _GEN_927;
  wire  _GEN_933 = 8'he8 == mshr_io_mshrInfo_index ? _T_257_232_1 : _GEN_929;
  wire  _GEN_934 = 8'he8 == mshr_io_mshrInfo_index ? _T_257_232_2 : _GEN_930;
  wire  _GEN_935 = 8'he8 == mshr_io_mshrInfo_index ? _T_257_232_3 : _GEN_931;
  wire  _GEN_937 = 8'he9 == mshr_io_mshrInfo_index ? _T_257_233_1 : _GEN_933;
  wire  _GEN_938 = 8'he9 == mshr_io_mshrInfo_index ? _T_257_233_2 : _GEN_934;
  wire  _GEN_939 = 8'he9 == mshr_io_mshrInfo_index ? _T_257_233_3 : _GEN_935;
  wire  _GEN_941 = 8'hea == mshr_io_mshrInfo_index ? _T_257_234_1 : _GEN_937;
  wire  _GEN_942 = 8'hea == mshr_io_mshrInfo_index ? _T_257_234_2 : _GEN_938;
  wire  _GEN_943 = 8'hea == mshr_io_mshrInfo_index ? _T_257_234_3 : _GEN_939;
  wire  _GEN_945 = 8'heb == mshr_io_mshrInfo_index ? _T_257_235_1 : _GEN_941;
  wire  _GEN_946 = 8'heb == mshr_io_mshrInfo_index ? _T_257_235_2 : _GEN_942;
  wire  _GEN_947 = 8'heb == mshr_io_mshrInfo_index ? _T_257_235_3 : _GEN_943;
  wire  _GEN_949 = 8'hec == mshr_io_mshrInfo_index ? _T_257_236_1 : _GEN_945;
  wire  _GEN_950 = 8'hec == mshr_io_mshrInfo_index ? _T_257_236_2 : _GEN_946;
  wire  _GEN_951 = 8'hec == mshr_io_mshrInfo_index ? _T_257_236_3 : _GEN_947;
  wire  _GEN_953 = 8'hed == mshr_io_mshrInfo_index ? _T_257_237_1 : _GEN_949;
  wire  _GEN_954 = 8'hed == mshr_io_mshrInfo_index ? _T_257_237_2 : _GEN_950;
  wire  _GEN_955 = 8'hed == mshr_io_mshrInfo_index ? _T_257_237_3 : _GEN_951;
  wire  _GEN_957 = 8'hee == mshr_io_mshrInfo_index ? _T_257_238_1 : _GEN_953;
  wire  _GEN_958 = 8'hee == mshr_io_mshrInfo_index ? _T_257_238_2 : _GEN_954;
  wire  _GEN_959 = 8'hee == mshr_io_mshrInfo_index ? _T_257_238_3 : _GEN_955;
  wire  _GEN_961 = 8'hef == mshr_io_mshrInfo_index ? _T_257_239_1 : _GEN_957;
  wire  _GEN_962 = 8'hef == mshr_io_mshrInfo_index ? _T_257_239_2 : _GEN_958;
  wire  _GEN_963 = 8'hef == mshr_io_mshrInfo_index ? _T_257_239_3 : _GEN_959;
  wire  _GEN_965 = 8'hf0 == mshr_io_mshrInfo_index ? _T_257_240_1 : _GEN_961;
  wire  _GEN_966 = 8'hf0 == mshr_io_mshrInfo_index ? _T_257_240_2 : _GEN_962;
  wire  _GEN_967 = 8'hf0 == mshr_io_mshrInfo_index ? _T_257_240_3 : _GEN_963;
  wire  _GEN_969 = 8'hf1 == mshr_io_mshrInfo_index ? _T_257_241_1 : _GEN_965;
  wire  _GEN_970 = 8'hf1 == mshr_io_mshrInfo_index ? _T_257_241_2 : _GEN_966;
  wire  _GEN_971 = 8'hf1 == mshr_io_mshrInfo_index ? _T_257_241_3 : _GEN_967;
  wire  _GEN_973 = 8'hf2 == mshr_io_mshrInfo_index ? _T_257_242_1 : _GEN_969;
  wire  _GEN_974 = 8'hf2 == mshr_io_mshrInfo_index ? _T_257_242_2 : _GEN_970;
  wire  _GEN_975 = 8'hf2 == mshr_io_mshrInfo_index ? _T_257_242_3 : _GEN_971;
  wire  _GEN_977 = 8'hf3 == mshr_io_mshrInfo_index ? _T_257_243_1 : _GEN_973;
  wire  _GEN_978 = 8'hf3 == mshr_io_mshrInfo_index ? _T_257_243_2 : _GEN_974;
  wire  _GEN_979 = 8'hf3 == mshr_io_mshrInfo_index ? _T_257_243_3 : _GEN_975;
  wire  _GEN_981 = 8'hf4 == mshr_io_mshrInfo_index ? _T_257_244_1 : _GEN_977;
  wire  _GEN_982 = 8'hf4 == mshr_io_mshrInfo_index ? _T_257_244_2 : _GEN_978;
  wire  _GEN_983 = 8'hf4 == mshr_io_mshrInfo_index ? _T_257_244_3 : _GEN_979;
  wire  _GEN_985 = 8'hf5 == mshr_io_mshrInfo_index ? _T_257_245_1 : _GEN_981;
  wire  _GEN_986 = 8'hf5 == mshr_io_mshrInfo_index ? _T_257_245_2 : _GEN_982;
  wire  _GEN_987 = 8'hf5 == mshr_io_mshrInfo_index ? _T_257_245_3 : _GEN_983;
  wire  _GEN_989 = 8'hf6 == mshr_io_mshrInfo_index ? _T_257_246_1 : _GEN_985;
  wire  _GEN_990 = 8'hf6 == mshr_io_mshrInfo_index ? _T_257_246_2 : _GEN_986;
  wire  _GEN_991 = 8'hf6 == mshr_io_mshrInfo_index ? _T_257_246_3 : _GEN_987;
  wire  _GEN_993 = 8'hf7 == mshr_io_mshrInfo_index ? _T_257_247_1 : _GEN_989;
  wire  _GEN_994 = 8'hf7 == mshr_io_mshrInfo_index ? _T_257_247_2 : _GEN_990;
  wire  _GEN_995 = 8'hf7 == mshr_io_mshrInfo_index ? _T_257_247_3 : _GEN_991;
  wire  _GEN_997 = 8'hf8 == mshr_io_mshrInfo_index ? _T_257_248_1 : _GEN_993;
  wire  _GEN_998 = 8'hf8 == mshr_io_mshrInfo_index ? _T_257_248_2 : _GEN_994;
  wire  _GEN_999 = 8'hf8 == mshr_io_mshrInfo_index ? _T_257_248_3 : _GEN_995;
  wire  _GEN_1001 = 8'hf9 == mshr_io_mshrInfo_index ? _T_257_249_1 : _GEN_997;
  wire  _GEN_1002 = 8'hf9 == mshr_io_mshrInfo_index ? _T_257_249_2 : _GEN_998;
  wire  _GEN_1003 = 8'hf9 == mshr_io_mshrInfo_index ? _T_257_249_3 : _GEN_999;
  wire  _GEN_1005 = 8'hfa == mshr_io_mshrInfo_index ? _T_257_250_1 : _GEN_1001;
  wire  _GEN_1006 = 8'hfa == mshr_io_mshrInfo_index ? _T_257_250_2 : _GEN_1002;
  wire  _GEN_1007 = 8'hfa == mshr_io_mshrInfo_index ? _T_257_250_3 : _GEN_1003;
  wire  _GEN_1009 = 8'hfb == mshr_io_mshrInfo_index ? _T_257_251_1 : _GEN_1005;
  wire  _GEN_1010 = 8'hfb == mshr_io_mshrInfo_index ? _T_257_251_2 : _GEN_1006;
  wire  _GEN_1011 = 8'hfb == mshr_io_mshrInfo_index ? _T_257_251_3 : _GEN_1007;
  wire  _GEN_1013 = 8'hfc == mshr_io_mshrInfo_index ? _T_257_252_1 : _GEN_1009;
  wire  _GEN_1014 = 8'hfc == mshr_io_mshrInfo_index ? _T_257_252_2 : _GEN_1010;
  wire  _GEN_1015 = 8'hfc == mshr_io_mshrInfo_index ? _T_257_252_3 : _GEN_1011;
  wire  _GEN_1017 = 8'hfd == mshr_io_mshrInfo_index ? _T_257_253_1 : _GEN_1013;
  wire  _GEN_1018 = 8'hfd == mshr_io_mshrInfo_index ? _T_257_253_2 : _GEN_1014;
  wire  _GEN_1019 = 8'hfd == mshr_io_mshrInfo_index ? _T_257_253_3 : _GEN_1015;
  wire  _GEN_1021 = 8'hfe == mshr_io_mshrInfo_index ? _T_257_254_1 : _GEN_1017;
  wire  _GEN_1022 = 8'hfe == mshr_io_mshrInfo_index ? _T_257_254_2 : _GEN_1018;
  wire  _GEN_1023 = 8'hfe == mshr_io_mshrInfo_index ? _T_257_254_3 : _GEN_1019;
  wire  _GEN_1025 = 8'hff == mshr_io_mshrInfo_index ? _T_257_255_1 : _GEN_1021;
  wire  _GEN_1026 = 8'hff == mshr_io_mshrInfo_index ? _T_257_255_2 : _GEN_1022;
  wire  _GEN_1027 = 8'hff == mshr_io_mshrInfo_index ? _T_257_255_3 : _GEN_1023;
  wire  _T_271 = ~_GEN_1025; // @[PLRUMRUNM.scala 42:43]
  wire  _T_272 = ~_GEN_1026; // @[PLRUMRUNM.scala 42:43]
  wire  _T_273 = ~_GEN_1027; // @[PLRUMRUNM.scala 42:43]
  wire [1:0] _T_275 = _T_272 ? 2'h2 : {{1'd0}, _T_271}; // @[PLRUMRUNM.scala 42:32]
  wire  _T_278 = ~io_data_ready; // @[QueryTop.scala 98:45]
  wire  _T_280 = ~readHolder_io_output_valid; // @[QueryTop.scala 103:42]
  wire  _T_281 = comparator_io_bankHitWay_valid & _T_280; // @[QueryTop.scala 103:39]
  wire [31:0] _T_282 = _T_281 ? _GEN_3 : readHolder_io_output_bits; // @[Mux.scala 98:16]
  wire [30:0] _T_286 = {io_fetchQuery_phyTag,io_fetchQuery_index,io_fetchQuery_bankIndex,2'h0}; // @[Cat.scala 29:58]
  wire [30:0] _T_289 = {mshr_io_mshrInfo_tag,mshr_io_mshrInfo_index,mshr_io_mshrInfo_bankIndex,2'h0}; // @[Cat.scala 29:58]
  wire [30:0] _T_290 = newMiss ? _T_286 : _T_289; // @[QueryTop.scala 107:29]
  wire  _T_291 = ~queryHit; // @[QueryTop.scala 120:38]
  wire  _GEN_1032 = 8'h1 == io_fetchQuery_index ? _T_257_1_0 : _T_257_0_0;
  wire  _GEN_1033 = 8'h1 == io_fetchQuery_index ? _T_257_1_1 : _T_257_0_1;
  wire  _GEN_1034 = 8'h1 == io_fetchQuery_index ? _T_257_1_2 : _T_257_0_2;
  wire  _GEN_1035 = 8'h1 == io_fetchQuery_index ? _T_257_1_3 : _T_257_0_3;
  wire  _GEN_1036 = 8'h2 == io_fetchQuery_index ? _T_257_2_0 : _GEN_1032;
  wire  _GEN_1037 = 8'h2 == io_fetchQuery_index ? _T_257_2_1 : _GEN_1033;
  wire  _GEN_1038 = 8'h2 == io_fetchQuery_index ? _T_257_2_2 : _GEN_1034;
  wire  _GEN_1039 = 8'h2 == io_fetchQuery_index ? _T_257_2_3 : _GEN_1035;
  wire  _GEN_1040 = 8'h3 == io_fetchQuery_index ? _T_257_3_0 : _GEN_1036;
  wire  _GEN_1041 = 8'h3 == io_fetchQuery_index ? _T_257_3_1 : _GEN_1037;
  wire  _GEN_1042 = 8'h3 == io_fetchQuery_index ? _T_257_3_2 : _GEN_1038;
  wire  _GEN_1043 = 8'h3 == io_fetchQuery_index ? _T_257_3_3 : _GEN_1039;
  wire  _GEN_1044 = 8'h4 == io_fetchQuery_index ? _T_257_4_0 : _GEN_1040;
  wire  _GEN_1045 = 8'h4 == io_fetchQuery_index ? _T_257_4_1 : _GEN_1041;
  wire  _GEN_1046 = 8'h4 == io_fetchQuery_index ? _T_257_4_2 : _GEN_1042;
  wire  _GEN_1047 = 8'h4 == io_fetchQuery_index ? _T_257_4_3 : _GEN_1043;
  wire  _GEN_1048 = 8'h5 == io_fetchQuery_index ? _T_257_5_0 : _GEN_1044;
  wire  _GEN_1049 = 8'h5 == io_fetchQuery_index ? _T_257_5_1 : _GEN_1045;
  wire  _GEN_1050 = 8'h5 == io_fetchQuery_index ? _T_257_5_2 : _GEN_1046;
  wire  _GEN_1051 = 8'h5 == io_fetchQuery_index ? _T_257_5_3 : _GEN_1047;
  wire  _GEN_1052 = 8'h6 == io_fetchQuery_index ? _T_257_6_0 : _GEN_1048;
  wire  _GEN_1053 = 8'h6 == io_fetchQuery_index ? _T_257_6_1 : _GEN_1049;
  wire  _GEN_1054 = 8'h6 == io_fetchQuery_index ? _T_257_6_2 : _GEN_1050;
  wire  _GEN_1055 = 8'h6 == io_fetchQuery_index ? _T_257_6_3 : _GEN_1051;
  wire  _GEN_1056 = 8'h7 == io_fetchQuery_index ? _T_257_7_0 : _GEN_1052;
  wire  _GEN_1057 = 8'h7 == io_fetchQuery_index ? _T_257_7_1 : _GEN_1053;
  wire  _GEN_1058 = 8'h7 == io_fetchQuery_index ? _T_257_7_2 : _GEN_1054;
  wire  _GEN_1059 = 8'h7 == io_fetchQuery_index ? _T_257_7_3 : _GEN_1055;
  wire  _GEN_1060 = 8'h8 == io_fetchQuery_index ? _T_257_8_0 : _GEN_1056;
  wire  _GEN_1061 = 8'h8 == io_fetchQuery_index ? _T_257_8_1 : _GEN_1057;
  wire  _GEN_1062 = 8'h8 == io_fetchQuery_index ? _T_257_8_2 : _GEN_1058;
  wire  _GEN_1063 = 8'h8 == io_fetchQuery_index ? _T_257_8_3 : _GEN_1059;
  wire  _GEN_1064 = 8'h9 == io_fetchQuery_index ? _T_257_9_0 : _GEN_1060;
  wire  _GEN_1065 = 8'h9 == io_fetchQuery_index ? _T_257_9_1 : _GEN_1061;
  wire  _GEN_1066 = 8'h9 == io_fetchQuery_index ? _T_257_9_2 : _GEN_1062;
  wire  _GEN_1067 = 8'h9 == io_fetchQuery_index ? _T_257_9_3 : _GEN_1063;
  wire  _GEN_1068 = 8'ha == io_fetchQuery_index ? _T_257_10_0 : _GEN_1064;
  wire  _GEN_1069 = 8'ha == io_fetchQuery_index ? _T_257_10_1 : _GEN_1065;
  wire  _GEN_1070 = 8'ha == io_fetchQuery_index ? _T_257_10_2 : _GEN_1066;
  wire  _GEN_1071 = 8'ha == io_fetchQuery_index ? _T_257_10_3 : _GEN_1067;
  wire  _GEN_1072 = 8'hb == io_fetchQuery_index ? _T_257_11_0 : _GEN_1068;
  wire  _GEN_1073 = 8'hb == io_fetchQuery_index ? _T_257_11_1 : _GEN_1069;
  wire  _GEN_1074 = 8'hb == io_fetchQuery_index ? _T_257_11_2 : _GEN_1070;
  wire  _GEN_1075 = 8'hb == io_fetchQuery_index ? _T_257_11_3 : _GEN_1071;
  wire  _GEN_1076 = 8'hc == io_fetchQuery_index ? _T_257_12_0 : _GEN_1072;
  wire  _GEN_1077 = 8'hc == io_fetchQuery_index ? _T_257_12_1 : _GEN_1073;
  wire  _GEN_1078 = 8'hc == io_fetchQuery_index ? _T_257_12_2 : _GEN_1074;
  wire  _GEN_1079 = 8'hc == io_fetchQuery_index ? _T_257_12_3 : _GEN_1075;
  wire  _GEN_1080 = 8'hd == io_fetchQuery_index ? _T_257_13_0 : _GEN_1076;
  wire  _GEN_1081 = 8'hd == io_fetchQuery_index ? _T_257_13_1 : _GEN_1077;
  wire  _GEN_1082 = 8'hd == io_fetchQuery_index ? _T_257_13_2 : _GEN_1078;
  wire  _GEN_1083 = 8'hd == io_fetchQuery_index ? _T_257_13_3 : _GEN_1079;
  wire  _GEN_1084 = 8'he == io_fetchQuery_index ? _T_257_14_0 : _GEN_1080;
  wire  _GEN_1085 = 8'he == io_fetchQuery_index ? _T_257_14_1 : _GEN_1081;
  wire  _GEN_1086 = 8'he == io_fetchQuery_index ? _T_257_14_2 : _GEN_1082;
  wire  _GEN_1087 = 8'he == io_fetchQuery_index ? _T_257_14_3 : _GEN_1083;
  wire  _GEN_1088 = 8'hf == io_fetchQuery_index ? _T_257_15_0 : _GEN_1084;
  wire  _GEN_1089 = 8'hf == io_fetchQuery_index ? _T_257_15_1 : _GEN_1085;
  wire  _GEN_1090 = 8'hf == io_fetchQuery_index ? _T_257_15_2 : _GEN_1086;
  wire  _GEN_1091 = 8'hf == io_fetchQuery_index ? _T_257_15_3 : _GEN_1087;
  wire  _GEN_1092 = 8'h10 == io_fetchQuery_index ? _T_257_16_0 : _GEN_1088;
  wire  _GEN_1093 = 8'h10 == io_fetchQuery_index ? _T_257_16_1 : _GEN_1089;
  wire  _GEN_1094 = 8'h10 == io_fetchQuery_index ? _T_257_16_2 : _GEN_1090;
  wire  _GEN_1095 = 8'h10 == io_fetchQuery_index ? _T_257_16_3 : _GEN_1091;
  wire  _GEN_1096 = 8'h11 == io_fetchQuery_index ? _T_257_17_0 : _GEN_1092;
  wire  _GEN_1097 = 8'h11 == io_fetchQuery_index ? _T_257_17_1 : _GEN_1093;
  wire  _GEN_1098 = 8'h11 == io_fetchQuery_index ? _T_257_17_2 : _GEN_1094;
  wire  _GEN_1099 = 8'h11 == io_fetchQuery_index ? _T_257_17_3 : _GEN_1095;
  wire  _GEN_1100 = 8'h12 == io_fetchQuery_index ? _T_257_18_0 : _GEN_1096;
  wire  _GEN_1101 = 8'h12 == io_fetchQuery_index ? _T_257_18_1 : _GEN_1097;
  wire  _GEN_1102 = 8'h12 == io_fetchQuery_index ? _T_257_18_2 : _GEN_1098;
  wire  _GEN_1103 = 8'h12 == io_fetchQuery_index ? _T_257_18_3 : _GEN_1099;
  wire  _GEN_1104 = 8'h13 == io_fetchQuery_index ? _T_257_19_0 : _GEN_1100;
  wire  _GEN_1105 = 8'h13 == io_fetchQuery_index ? _T_257_19_1 : _GEN_1101;
  wire  _GEN_1106 = 8'h13 == io_fetchQuery_index ? _T_257_19_2 : _GEN_1102;
  wire  _GEN_1107 = 8'h13 == io_fetchQuery_index ? _T_257_19_3 : _GEN_1103;
  wire  _GEN_1108 = 8'h14 == io_fetchQuery_index ? _T_257_20_0 : _GEN_1104;
  wire  _GEN_1109 = 8'h14 == io_fetchQuery_index ? _T_257_20_1 : _GEN_1105;
  wire  _GEN_1110 = 8'h14 == io_fetchQuery_index ? _T_257_20_2 : _GEN_1106;
  wire  _GEN_1111 = 8'h14 == io_fetchQuery_index ? _T_257_20_3 : _GEN_1107;
  wire  _GEN_1112 = 8'h15 == io_fetchQuery_index ? _T_257_21_0 : _GEN_1108;
  wire  _GEN_1113 = 8'h15 == io_fetchQuery_index ? _T_257_21_1 : _GEN_1109;
  wire  _GEN_1114 = 8'h15 == io_fetchQuery_index ? _T_257_21_2 : _GEN_1110;
  wire  _GEN_1115 = 8'h15 == io_fetchQuery_index ? _T_257_21_3 : _GEN_1111;
  wire  _GEN_1116 = 8'h16 == io_fetchQuery_index ? _T_257_22_0 : _GEN_1112;
  wire  _GEN_1117 = 8'h16 == io_fetchQuery_index ? _T_257_22_1 : _GEN_1113;
  wire  _GEN_1118 = 8'h16 == io_fetchQuery_index ? _T_257_22_2 : _GEN_1114;
  wire  _GEN_1119 = 8'h16 == io_fetchQuery_index ? _T_257_22_3 : _GEN_1115;
  wire  _GEN_1120 = 8'h17 == io_fetchQuery_index ? _T_257_23_0 : _GEN_1116;
  wire  _GEN_1121 = 8'h17 == io_fetchQuery_index ? _T_257_23_1 : _GEN_1117;
  wire  _GEN_1122 = 8'h17 == io_fetchQuery_index ? _T_257_23_2 : _GEN_1118;
  wire  _GEN_1123 = 8'h17 == io_fetchQuery_index ? _T_257_23_3 : _GEN_1119;
  wire  _GEN_1124 = 8'h18 == io_fetchQuery_index ? _T_257_24_0 : _GEN_1120;
  wire  _GEN_1125 = 8'h18 == io_fetchQuery_index ? _T_257_24_1 : _GEN_1121;
  wire  _GEN_1126 = 8'h18 == io_fetchQuery_index ? _T_257_24_2 : _GEN_1122;
  wire  _GEN_1127 = 8'h18 == io_fetchQuery_index ? _T_257_24_3 : _GEN_1123;
  wire  _GEN_1128 = 8'h19 == io_fetchQuery_index ? _T_257_25_0 : _GEN_1124;
  wire  _GEN_1129 = 8'h19 == io_fetchQuery_index ? _T_257_25_1 : _GEN_1125;
  wire  _GEN_1130 = 8'h19 == io_fetchQuery_index ? _T_257_25_2 : _GEN_1126;
  wire  _GEN_1131 = 8'h19 == io_fetchQuery_index ? _T_257_25_3 : _GEN_1127;
  wire  _GEN_1132 = 8'h1a == io_fetchQuery_index ? _T_257_26_0 : _GEN_1128;
  wire  _GEN_1133 = 8'h1a == io_fetchQuery_index ? _T_257_26_1 : _GEN_1129;
  wire  _GEN_1134 = 8'h1a == io_fetchQuery_index ? _T_257_26_2 : _GEN_1130;
  wire  _GEN_1135 = 8'h1a == io_fetchQuery_index ? _T_257_26_3 : _GEN_1131;
  wire  _GEN_1136 = 8'h1b == io_fetchQuery_index ? _T_257_27_0 : _GEN_1132;
  wire  _GEN_1137 = 8'h1b == io_fetchQuery_index ? _T_257_27_1 : _GEN_1133;
  wire  _GEN_1138 = 8'h1b == io_fetchQuery_index ? _T_257_27_2 : _GEN_1134;
  wire  _GEN_1139 = 8'h1b == io_fetchQuery_index ? _T_257_27_3 : _GEN_1135;
  wire  _GEN_1140 = 8'h1c == io_fetchQuery_index ? _T_257_28_0 : _GEN_1136;
  wire  _GEN_1141 = 8'h1c == io_fetchQuery_index ? _T_257_28_1 : _GEN_1137;
  wire  _GEN_1142 = 8'h1c == io_fetchQuery_index ? _T_257_28_2 : _GEN_1138;
  wire  _GEN_1143 = 8'h1c == io_fetchQuery_index ? _T_257_28_3 : _GEN_1139;
  wire  _GEN_1144 = 8'h1d == io_fetchQuery_index ? _T_257_29_0 : _GEN_1140;
  wire  _GEN_1145 = 8'h1d == io_fetchQuery_index ? _T_257_29_1 : _GEN_1141;
  wire  _GEN_1146 = 8'h1d == io_fetchQuery_index ? _T_257_29_2 : _GEN_1142;
  wire  _GEN_1147 = 8'h1d == io_fetchQuery_index ? _T_257_29_3 : _GEN_1143;
  wire  _GEN_1148 = 8'h1e == io_fetchQuery_index ? _T_257_30_0 : _GEN_1144;
  wire  _GEN_1149 = 8'h1e == io_fetchQuery_index ? _T_257_30_1 : _GEN_1145;
  wire  _GEN_1150 = 8'h1e == io_fetchQuery_index ? _T_257_30_2 : _GEN_1146;
  wire  _GEN_1151 = 8'h1e == io_fetchQuery_index ? _T_257_30_3 : _GEN_1147;
  wire  _GEN_1152 = 8'h1f == io_fetchQuery_index ? _T_257_31_0 : _GEN_1148;
  wire  _GEN_1153 = 8'h1f == io_fetchQuery_index ? _T_257_31_1 : _GEN_1149;
  wire  _GEN_1154 = 8'h1f == io_fetchQuery_index ? _T_257_31_2 : _GEN_1150;
  wire  _GEN_1155 = 8'h1f == io_fetchQuery_index ? _T_257_31_3 : _GEN_1151;
  wire  _GEN_1156 = 8'h20 == io_fetchQuery_index ? _T_257_32_0 : _GEN_1152;
  wire  _GEN_1157 = 8'h20 == io_fetchQuery_index ? _T_257_32_1 : _GEN_1153;
  wire  _GEN_1158 = 8'h20 == io_fetchQuery_index ? _T_257_32_2 : _GEN_1154;
  wire  _GEN_1159 = 8'h20 == io_fetchQuery_index ? _T_257_32_3 : _GEN_1155;
  wire  _GEN_1160 = 8'h21 == io_fetchQuery_index ? _T_257_33_0 : _GEN_1156;
  wire  _GEN_1161 = 8'h21 == io_fetchQuery_index ? _T_257_33_1 : _GEN_1157;
  wire  _GEN_1162 = 8'h21 == io_fetchQuery_index ? _T_257_33_2 : _GEN_1158;
  wire  _GEN_1163 = 8'h21 == io_fetchQuery_index ? _T_257_33_3 : _GEN_1159;
  wire  _GEN_1164 = 8'h22 == io_fetchQuery_index ? _T_257_34_0 : _GEN_1160;
  wire  _GEN_1165 = 8'h22 == io_fetchQuery_index ? _T_257_34_1 : _GEN_1161;
  wire  _GEN_1166 = 8'h22 == io_fetchQuery_index ? _T_257_34_2 : _GEN_1162;
  wire  _GEN_1167 = 8'h22 == io_fetchQuery_index ? _T_257_34_3 : _GEN_1163;
  wire  _GEN_1168 = 8'h23 == io_fetchQuery_index ? _T_257_35_0 : _GEN_1164;
  wire  _GEN_1169 = 8'h23 == io_fetchQuery_index ? _T_257_35_1 : _GEN_1165;
  wire  _GEN_1170 = 8'h23 == io_fetchQuery_index ? _T_257_35_2 : _GEN_1166;
  wire  _GEN_1171 = 8'h23 == io_fetchQuery_index ? _T_257_35_3 : _GEN_1167;
  wire  _GEN_1172 = 8'h24 == io_fetchQuery_index ? _T_257_36_0 : _GEN_1168;
  wire  _GEN_1173 = 8'h24 == io_fetchQuery_index ? _T_257_36_1 : _GEN_1169;
  wire  _GEN_1174 = 8'h24 == io_fetchQuery_index ? _T_257_36_2 : _GEN_1170;
  wire  _GEN_1175 = 8'h24 == io_fetchQuery_index ? _T_257_36_3 : _GEN_1171;
  wire  _GEN_1176 = 8'h25 == io_fetchQuery_index ? _T_257_37_0 : _GEN_1172;
  wire  _GEN_1177 = 8'h25 == io_fetchQuery_index ? _T_257_37_1 : _GEN_1173;
  wire  _GEN_1178 = 8'h25 == io_fetchQuery_index ? _T_257_37_2 : _GEN_1174;
  wire  _GEN_1179 = 8'h25 == io_fetchQuery_index ? _T_257_37_3 : _GEN_1175;
  wire  _GEN_1180 = 8'h26 == io_fetchQuery_index ? _T_257_38_0 : _GEN_1176;
  wire  _GEN_1181 = 8'h26 == io_fetchQuery_index ? _T_257_38_1 : _GEN_1177;
  wire  _GEN_1182 = 8'h26 == io_fetchQuery_index ? _T_257_38_2 : _GEN_1178;
  wire  _GEN_1183 = 8'h26 == io_fetchQuery_index ? _T_257_38_3 : _GEN_1179;
  wire  _GEN_1184 = 8'h27 == io_fetchQuery_index ? _T_257_39_0 : _GEN_1180;
  wire  _GEN_1185 = 8'h27 == io_fetchQuery_index ? _T_257_39_1 : _GEN_1181;
  wire  _GEN_1186 = 8'h27 == io_fetchQuery_index ? _T_257_39_2 : _GEN_1182;
  wire  _GEN_1187 = 8'h27 == io_fetchQuery_index ? _T_257_39_3 : _GEN_1183;
  wire  _GEN_1188 = 8'h28 == io_fetchQuery_index ? _T_257_40_0 : _GEN_1184;
  wire  _GEN_1189 = 8'h28 == io_fetchQuery_index ? _T_257_40_1 : _GEN_1185;
  wire  _GEN_1190 = 8'h28 == io_fetchQuery_index ? _T_257_40_2 : _GEN_1186;
  wire  _GEN_1191 = 8'h28 == io_fetchQuery_index ? _T_257_40_3 : _GEN_1187;
  wire  _GEN_1192 = 8'h29 == io_fetchQuery_index ? _T_257_41_0 : _GEN_1188;
  wire  _GEN_1193 = 8'h29 == io_fetchQuery_index ? _T_257_41_1 : _GEN_1189;
  wire  _GEN_1194 = 8'h29 == io_fetchQuery_index ? _T_257_41_2 : _GEN_1190;
  wire  _GEN_1195 = 8'h29 == io_fetchQuery_index ? _T_257_41_3 : _GEN_1191;
  wire  _GEN_1196 = 8'h2a == io_fetchQuery_index ? _T_257_42_0 : _GEN_1192;
  wire  _GEN_1197 = 8'h2a == io_fetchQuery_index ? _T_257_42_1 : _GEN_1193;
  wire  _GEN_1198 = 8'h2a == io_fetchQuery_index ? _T_257_42_2 : _GEN_1194;
  wire  _GEN_1199 = 8'h2a == io_fetchQuery_index ? _T_257_42_3 : _GEN_1195;
  wire  _GEN_1200 = 8'h2b == io_fetchQuery_index ? _T_257_43_0 : _GEN_1196;
  wire  _GEN_1201 = 8'h2b == io_fetchQuery_index ? _T_257_43_1 : _GEN_1197;
  wire  _GEN_1202 = 8'h2b == io_fetchQuery_index ? _T_257_43_2 : _GEN_1198;
  wire  _GEN_1203 = 8'h2b == io_fetchQuery_index ? _T_257_43_3 : _GEN_1199;
  wire  _GEN_1204 = 8'h2c == io_fetchQuery_index ? _T_257_44_0 : _GEN_1200;
  wire  _GEN_1205 = 8'h2c == io_fetchQuery_index ? _T_257_44_1 : _GEN_1201;
  wire  _GEN_1206 = 8'h2c == io_fetchQuery_index ? _T_257_44_2 : _GEN_1202;
  wire  _GEN_1207 = 8'h2c == io_fetchQuery_index ? _T_257_44_3 : _GEN_1203;
  wire  _GEN_1208 = 8'h2d == io_fetchQuery_index ? _T_257_45_0 : _GEN_1204;
  wire  _GEN_1209 = 8'h2d == io_fetchQuery_index ? _T_257_45_1 : _GEN_1205;
  wire  _GEN_1210 = 8'h2d == io_fetchQuery_index ? _T_257_45_2 : _GEN_1206;
  wire  _GEN_1211 = 8'h2d == io_fetchQuery_index ? _T_257_45_3 : _GEN_1207;
  wire  _GEN_1212 = 8'h2e == io_fetchQuery_index ? _T_257_46_0 : _GEN_1208;
  wire  _GEN_1213 = 8'h2e == io_fetchQuery_index ? _T_257_46_1 : _GEN_1209;
  wire  _GEN_1214 = 8'h2e == io_fetchQuery_index ? _T_257_46_2 : _GEN_1210;
  wire  _GEN_1215 = 8'h2e == io_fetchQuery_index ? _T_257_46_3 : _GEN_1211;
  wire  _GEN_1216 = 8'h2f == io_fetchQuery_index ? _T_257_47_0 : _GEN_1212;
  wire  _GEN_1217 = 8'h2f == io_fetchQuery_index ? _T_257_47_1 : _GEN_1213;
  wire  _GEN_1218 = 8'h2f == io_fetchQuery_index ? _T_257_47_2 : _GEN_1214;
  wire  _GEN_1219 = 8'h2f == io_fetchQuery_index ? _T_257_47_3 : _GEN_1215;
  wire  _GEN_1220 = 8'h30 == io_fetchQuery_index ? _T_257_48_0 : _GEN_1216;
  wire  _GEN_1221 = 8'h30 == io_fetchQuery_index ? _T_257_48_1 : _GEN_1217;
  wire  _GEN_1222 = 8'h30 == io_fetchQuery_index ? _T_257_48_2 : _GEN_1218;
  wire  _GEN_1223 = 8'h30 == io_fetchQuery_index ? _T_257_48_3 : _GEN_1219;
  wire  _GEN_1224 = 8'h31 == io_fetchQuery_index ? _T_257_49_0 : _GEN_1220;
  wire  _GEN_1225 = 8'h31 == io_fetchQuery_index ? _T_257_49_1 : _GEN_1221;
  wire  _GEN_1226 = 8'h31 == io_fetchQuery_index ? _T_257_49_2 : _GEN_1222;
  wire  _GEN_1227 = 8'h31 == io_fetchQuery_index ? _T_257_49_3 : _GEN_1223;
  wire  _GEN_1228 = 8'h32 == io_fetchQuery_index ? _T_257_50_0 : _GEN_1224;
  wire  _GEN_1229 = 8'h32 == io_fetchQuery_index ? _T_257_50_1 : _GEN_1225;
  wire  _GEN_1230 = 8'h32 == io_fetchQuery_index ? _T_257_50_2 : _GEN_1226;
  wire  _GEN_1231 = 8'h32 == io_fetchQuery_index ? _T_257_50_3 : _GEN_1227;
  wire  _GEN_1232 = 8'h33 == io_fetchQuery_index ? _T_257_51_0 : _GEN_1228;
  wire  _GEN_1233 = 8'h33 == io_fetchQuery_index ? _T_257_51_1 : _GEN_1229;
  wire  _GEN_1234 = 8'h33 == io_fetchQuery_index ? _T_257_51_2 : _GEN_1230;
  wire  _GEN_1235 = 8'h33 == io_fetchQuery_index ? _T_257_51_3 : _GEN_1231;
  wire  _GEN_1236 = 8'h34 == io_fetchQuery_index ? _T_257_52_0 : _GEN_1232;
  wire  _GEN_1237 = 8'h34 == io_fetchQuery_index ? _T_257_52_1 : _GEN_1233;
  wire  _GEN_1238 = 8'h34 == io_fetchQuery_index ? _T_257_52_2 : _GEN_1234;
  wire  _GEN_1239 = 8'h34 == io_fetchQuery_index ? _T_257_52_3 : _GEN_1235;
  wire  _GEN_1240 = 8'h35 == io_fetchQuery_index ? _T_257_53_0 : _GEN_1236;
  wire  _GEN_1241 = 8'h35 == io_fetchQuery_index ? _T_257_53_1 : _GEN_1237;
  wire  _GEN_1242 = 8'h35 == io_fetchQuery_index ? _T_257_53_2 : _GEN_1238;
  wire  _GEN_1243 = 8'h35 == io_fetchQuery_index ? _T_257_53_3 : _GEN_1239;
  wire  _GEN_1244 = 8'h36 == io_fetchQuery_index ? _T_257_54_0 : _GEN_1240;
  wire  _GEN_1245 = 8'h36 == io_fetchQuery_index ? _T_257_54_1 : _GEN_1241;
  wire  _GEN_1246 = 8'h36 == io_fetchQuery_index ? _T_257_54_2 : _GEN_1242;
  wire  _GEN_1247 = 8'h36 == io_fetchQuery_index ? _T_257_54_3 : _GEN_1243;
  wire  _GEN_1248 = 8'h37 == io_fetchQuery_index ? _T_257_55_0 : _GEN_1244;
  wire  _GEN_1249 = 8'h37 == io_fetchQuery_index ? _T_257_55_1 : _GEN_1245;
  wire  _GEN_1250 = 8'h37 == io_fetchQuery_index ? _T_257_55_2 : _GEN_1246;
  wire  _GEN_1251 = 8'h37 == io_fetchQuery_index ? _T_257_55_3 : _GEN_1247;
  wire  _GEN_1252 = 8'h38 == io_fetchQuery_index ? _T_257_56_0 : _GEN_1248;
  wire  _GEN_1253 = 8'h38 == io_fetchQuery_index ? _T_257_56_1 : _GEN_1249;
  wire  _GEN_1254 = 8'h38 == io_fetchQuery_index ? _T_257_56_2 : _GEN_1250;
  wire  _GEN_1255 = 8'h38 == io_fetchQuery_index ? _T_257_56_3 : _GEN_1251;
  wire  _GEN_1256 = 8'h39 == io_fetchQuery_index ? _T_257_57_0 : _GEN_1252;
  wire  _GEN_1257 = 8'h39 == io_fetchQuery_index ? _T_257_57_1 : _GEN_1253;
  wire  _GEN_1258 = 8'h39 == io_fetchQuery_index ? _T_257_57_2 : _GEN_1254;
  wire  _GEN_1259 = 8'h39 == io_fetchQuery_index ? _T_257_57_3 : _GEN_1255;
  wire  _GEN_1260 = 8'h3a == io_fetchQuery_index ? _T_257_58_0 : _GEN_1256;
  wire  _GEN_1261 = 8'h3a == io_fetchQuery_index ? _T_257_58_1 : _GEN_1257;
  wire  _GEN_1262 = 8'h3a == io_fetchQuery_index ? _T_257_58_2 : _GEN_1258;
  wire  _GEN_1263 = 8'h3a == io_fetchQuery_index ? _T_257_58_3 : _GEN_1259;
  wire  _GEN_1264 = 8'h3b == io_fetchQuery_index ? _T_257_59_0 : _GEN_1260;
  wire  _GEN_1265 = 8'h3b == io_fetchQuery_index ? _T_257_59_1 : _GEN_1261;
  wire  _GEN_1266 = 8'h3b == io_fetchQuery_index ? _T_257_59_2 : _GEN_1262;
  wire  _GEN_1267 = 8'h3b == io_fetchQuery_index ? _T_257_59_3 : _GEN_1263;
  wire  _GEN_1268 = 8'h3c == io_fetchQuery_index ? _T_257_60_0 : _GEN_1264;
  wire  _GEN_1269 = 8'h3c == io_fetchQuery_index ? _T_257_60_1 : _GEN_1265;
  wire  _GEN_1270 = 8'h3c == io_fetchQuery_index ? _T_257_60_2 : _GEN_1266;
  wire  _GEN_1271 = 8'h3c == io_fetchQuery_index ? _T_257_60_3 : _GEN_1267;
  wire  _GEN_1272 = 8'h3d == io_fetchQuery_index ? _T_257_61_0 : _GEN_1268;
  wire  _GEN_1273 = 8'h3d == io_fetchQuery_index ? _T_257_61_1 : _GEN_1269;
  wire  _GEN_1274 = 8'h3d == io_fetchQuery_index ? _T_257_61_2 : _GEN_1270;
  wire  _GEN_1275 = 8'h3d == io_fetchQuery_index ? _T_257_61_3 : _GEN_1271;
  wire  _GEN_1276 = 8'h3e == io_fetchQuery_index ? _T_257_62_0 : _GEN_1272;
  wire  _GEN_1277 = 8'h3e == io_fetchQuery_index ? _T_257_62_1 : _GEN_1273;
  wire  _GEN_1278 = 8'h3e == io_fetchQuery_index ? _T_257_62_2 : _GEN_1274;
  wire  _GEN_1279 = 8'h3e == io_fetchQuery_index ? _T_257_62_3 : _GEN_1275;
  wire  _GEN_1280 = 8'h3f == io_fetchQuery_index ? _T_257_63_0 : _GEN_1276;
  wire  _GEN_1281 = 8'h3f == io_fetchQuery_index ? _T_257_63_1 : _GEN_1277;
  wire  _GEN_1282 = 8'h3f == io_fetchQuery_index ? _T_257_63_2 : _GEN_1278;
  wire  _GEN_1283 = 8'h3f == io_fetchQuery_index ? _T_257_63_3 : _GEN_1279;
  wire  _GEN_1284 = 8'h40 == io_fetchQuery_index ? _T_257_64_0 : _GEN_1280;
  wire  _GEN_1285 = 8'h40 == io_fetchQuery_index ? _T_257_64_1 : _GEN_1281;
  wire  _GEN_1286 = 8'h40 == io_fetchQuery_index ? _T_257_64_2 : _GEN_1282;
  wire  _GEN_1287 = 8'h40 == io_fetchQuery_index ? _T_257_64_3 : _GEN_1283;
  wire  _GEN_1288 = 8'h41 == io_fetchQuery_index ? _T_257_65_0 : _GEN_1284;
  wire  _GEN_1289 = 8'h41 == io_fetchQuery_index ? _T_257_65_1 : _GEN_1285;
  wire  _GEN_1290 = 8'h41 == io_fetchQuery_index ? _T_257_65_2 : _GEN_1286;
  wire  _GEN_1291 = 8'h41 == io_fetchQuery_index ? _T_257_65_3 : _GEN_1287;
  wire  _GEN_1292 = 8'h42 == io_fetchQuery_index ? _T_257_66_0 : _GEN_1288;
  wire  _GEN_1293 = 8'h42 == io_fetchQuery_index ? _T_257_66_1 : _GEN_1289;
  wire  _GEN_1294 = 8'h42 == io_fetchQuery_index ? _T_257_66_2 : _GEN_1290;
  wire  _GEN_1295 = 8'h42 == io_fetchQuery_index ? _T_257_66_3 : _GEN_1291;
  wire  _GEN_1296 = 8'h43 == io_fetchQuery_index ? _T_257_67_0 : _GEN_1292;
  wire  _GEN_1297 = 8'h43 == io_fetchQuery_index ? _T_257_67_1 : _GEN_1293;
  wire  _GEN_1298 = 8'h43 == io_fetchQuery_index ? _T_257_67_2 : _GEN_1294;
  wire  _GEN_1299 = 8'h43 == io_fetchQuery_index ? _T_257_67_3 : _GEN_1295;
  wire  _GEN_1300 = 8'h44 == io_fetchQuery_index ? _T_257_68_0 : _GEN_1296;
  wire  _GEN_1301 = 8'h44 == io_fetchQuery_index ? _T_257_68_1 : _GEN_1297;
  wire  _GEN_1302 = 8'h44 == io_fetchQuery_index ? _T_257_68_2 : _GEN_1298;
  wire  _GEN_1303 = 8'h44 == io_fetchQuery_index ? _T_257_68_3 : _GEN_1299;
  wire  _GEN_1304 = 8'h45 == io_fetchQuery_index ? _T_257_69_0 : _GEN_1300;
  wire  _GEN_1305 = 8'h45 == io_fetchQuery_index ? _T_257_69_1 : _GEN_1301;
  wire  _GEN_1306 = 8'h45 == io_fetchQuery_index ? _T_257_69_2 : _GEN_1302;
  wire  _GEN_1307 = 8'h45 == io_fetchQuery_index ? _T_257_69_3 : _GEN_1303;
  wire  _GEN_1308 = 8'h46 == io_fetchQuery_index ? _T_257_70_0 : _GEN_1304;
  wire  _GEN_1309 = 8'h46 == io_fetchQuery_index ? _T_257_70_1 : _GEN_1305;
  wire  _GEN_1310 = 8'h46 == io_fetchQuery_index ? _T_257_70_2 : _GEN_1306;
  wire  _GEN_1311 = 8'h46 == io_fetchQuery_index ? _T_257_70_3 : _GEN_1307;
  wire  _GEN_1312 = 8'h47 == io_fetchQuery_index ? _T_257_71_0 : _GEN_1308;
  wire  _GEN_1313 = 8'h47 == io_fetchQuery_index ? _T_257_71_1 : _GEN_1309;
  wire  _GEN_1314 = 8'h47 == io_fetchQuery_index ? _T_257_71_2 : _GEN_1310;
  wire  _GEN_1315 = 8'h47 == io_fetchQuery_index ? _T_257_71_3 : _GEN_1311;
  wire  _GEN_1316 = 8'h48 == io_fetchQuery_index ? _T_257_72_0 : _GEN_1312;
  wire  _GEN_1317 = 8'h48 == io_fetchQuery_index ? _T_257_72_1 : _GEN_1313;
  wire  _GEN_1318 = 8'h48 == io_fetchQuery_index ? _T_257_72_2 : _GEN_1314;
  wire  _GEN_1319 = 8'h48 == io_fetchQuery_index ? _T_257_72_3 : _GEN_1315;
  wire  _GEN_1320 = 8'h49 == io_fetchQuery_index ? _T_257_73_0 : _GEN_1316;
  wire  _GEN_1321 = 8'h49 == io_fetchQuery_index ? _T_257_73_1 : _GEN_1317;
  wire  _GEN_1322 = 8'h49 == io_fetchQuery_index ? _T_257_73_2 : _GEN_1318;
  wire  _GEN_1323 = 8'h49 == io_fetchQuery_index ? _T_257_73_3 : _GEN_1319;
  wire  _GEN_1324 = 8'h4a == io_fetchQuery_index ? _T_257_74_0 : _GEN_1320;
  wire  _GEN_1325 = 8'h4a == io_fetchQuery_index ? _T_257_74_1 : _GEN_1321;
  wire  _GEN_1326 = 8'h4a == io_fetchQuery_index ? _T_257_74_2 : _GEN_1322;
  wire  _GEN_1327 = 8'h4a == io_fetchQuery_index ? _T_257_74_3 : _GEN_1323;
  wire  _GEN_1328 = 8'h4b == io_fetchQuery_index ? _T_257_75_0 : _GEN_1324;
  wire  _GEN_1329 = 8'h4b == io_fetchQuery_index ? _T_257_75_1 : _GEN_1325;
  wire  _GEN_1330 = 8'h4b == io_fetchQuery_index ? _T_257_75_2 : _GEN_1326;
  wire  _GEN_1331 = 8'h4b == io_fetchQuery_index ? _T_257_75_3 : _GEN_1327;
  wire  _GEN_1332 = 8'h4c == io_fetchQuery_index ? _T_257_76_0 : _GEN_1328;
  wire  _GEN_1333 = 8'h4c == io_fetchQuery_index ? _T_257_76_1 : _GEN_1329;
  wire  _GEN_1334 = 8'h4c == io_fetchQuery_index ? _T_257_76_2 : _GEN_1330;
  wire  _GEN_1335 = 8'h4c == io_fetchQuery_index ? _T_257_76_3 : _GEN_1331;
  wire  _GEN_1336 = 8'h4d == io_fetchQuery_index ? _T_257_77_0 : _GEN_1332;
  wire  _GEN_1337 = 8'h4d == io_fetchQuery_index ? _T_257_77_1 : _GEN_1333;
  wire  _GEN_1338 = 8'h4d == io_fetchQuery_index ? _T_257_77_2 : _GEN_1334;
  wire  _GEN_1339 = 8'h4d == io_fetchQuery_index ? _T_257_77_3 : _GEN_1335;
  wire  _GEN_1340 = 8'h4e == io_fetchQuery_index ? _T_257_78_0 : _GEN_1336;
  wire  _GEN_1341 = 8'h4e == io_fetchQuery_index ? _T_257_78_1 : _GEN_1337;
  wire  _GEN_1342 = 8'h4e == io_fetchQuery_index ? _T_257_78_2 : _GEN_1338;
  wire  _GEN_1343 = 8'h4e == io_fetchQuery_index ? _T_257_78_3 : _GEN_1339;
  wire  _GEN_1344 = 8'h4f == io_fetchQuery_index ? _T_257_79_0 : _GEN_1340;
  wire  _GEN_1345 = 8'h4f == io_fetchQuery_index ? _T_257_79_1 : _GEN_1341;
  wire  _GEN_1346 = 8'h4f == io_fetchQuery_index ? _T_257_79_2 : _GEN_1342;
  wire  _GEN_1347 = 8'h4f == io_fetchQuery_index ? _T_257_79_3 : _GEN_1343;
  wire  _GEN_1348 = 8'h50 == io_fetchQuery_index ? _T_257_80_0 : _GEN_1344;
  wire  _GEN_1349 = 8'h50 == io_fetchQuery_index ? _T_257_80_1 : _GEN_1345;
  wire  _GEN_1350 = 8'h50 == io_fetchQuery_index ? _T_257_80_2 : _GEN_1346;
  wire  _GEN_1351 = 8'h50 == io_fetchQuery_index ? _T_257_80_3 : _GEN_1347;
  wire  _GEN_1352 = 8'h51 == io_fetchQuery_index ? _T_257_81_0 : _GEN_1348;
  wire  _GEN_1353 = 8'h51 == io_fetchQuery_index ? _T_257_81_1 : _GEN_1349;
  wire  _GEN_1354 = 8'h51 == io_fetchQuery_index ? _T_257_81_2 : _GEN_1350;
  wire  _GEN_1355 = 8'h51 == io_fetchQuery_index ? _T_257_81_3 : _GEN_1351;
  wire  _GEN_1356 = 8'h52 == io_fetchQuery_index ? _T_257_82_0 : _GEN_1352;
  wire  _GEN_1357 = 8'h52 == io_fetchQuery_index ? _T_257_82_1 : _GEN_1353;
  wire  _GEN_1358 = 8'h52 == io_fetchQuery_index ? _T_257_82_2 : _GEN_1354;
  wire  _GEN_1359 = 8'h52 == io_fetchQuery_index ? _T_257_82_3 : _GEN_1355;
  wire  _GEN_1360 = 8'h53 == io_fetchQuery_index ? _T_257_83_0 : _GEN_1356;
  wire  _GEN_1361 = 8'h53 == io_fetchQuery_index ? _T_257_83_1 : _GEN_1357;
  wire  _GEN_1362 = 8'h53 == io_fetchQuery_index ? _T_257_83_2 : _GEN_1358;
  wire  _GEN_1363 = 8'h53 == io_fetchQuery_index ? _T_257_83_3 : _GEN_1359;
  wire  _GEN_1364 = 8'h54 == io_fetchQuery_index ? _T_257_84_0 : _GEN_1360;
  wire  _GEN_1365 = 8'h54 == io_fetchQuery_index ? _T_257_84_1 : _GEN_1361;
  wire  _GEN_1366 = 8'h54 == io_fetchQuery_index ? _T_257_84_2 : _GEN_1362;
  wire  _GEN_1367 = 8'h54 == io_fetchQuery_index ? _T_257_84_3 : _GEN_1363;
  wire  _GEN_1368 = 8'h55 == io_fetchQuery_index ? _T_257_85_0 : _GEN_1364;
  wire  _GEN_1369 = 8'h55 == io_fetchQuery_index ? _T_257_85_1 : _GEN_1365;
  wire  _GEN_1370 = 8'h55 == io_fetchQuery_index ? _T_257_85_2 : _GEN_1366;
  wire  _GEN_1371 = 8'h55 == io_fetchQuery_index ? _T_257_85_3 : _GEN_1367;
  wire  _GEN_1372 = 8'h56 == io_fetchQuery_index ? _T_257_86_0 : _GEN_1368;
  wire  _GEN_1373 = 8'h56 == io_fetchQuery_index ? _T_257_86_1 : _GEN_1369;
  wire  _GEN_1374 = 8'h56 == io_fetchQuery_index ? _T_257_86_2 : _GEN_1370;
  wire  _GEN_1375 = 8'h56 == io_fetchQuery_index ? _T_257_86_3 : _GEN_1371;
  wire  _GEN_1376 = 8'h57 == io_fetchQuery_index ? _T_257_87_0 : _GEN_1372;
  wire  _GEN_1377 = 8'h57 == io_fetchQuery_index ? _T_257_87_1 : _GEN_1373;
  wire  _GEN_1378 = 8'h57 == io_fetchQuery_index ? _T_257_87_2 : _GEN_1374;
  wire  _GEN_1379 = 8'h57 == io_fetchQuery_index ? _T_257_87_3 : _GEN_1375;
  wire  _GEN_1380 = 8'h58 == io_fetchQuery_index ? _T_257_88_0 : _GEN_1376;
  wire  _GEN_1381 = 8'h58 == io_fetchQuery_index ? _T_257_88_1 : _GEN_1377;
  wire  _GEN_1382 = 8'h58 == io_fetchQuery_index ? _T_257_88_2 : _GEN_1378;
  wire  _GEN_1383 = 8'h58 == io_fetchQuery_index ? _T_257_88_3 : _GEN_1379;
  wire  _GEN_1384 = 8'h59 == io_fetchQuery_index ? _T_257_89_0 : _GEN_1380;
  wire  _GEN_1385 = 8'h59 == io_fetchQuery_index ? _T_257_89_1 : _GEN_1381;
  wire  _GEN_1386 = 8'h59 == io_fetchQuery_index ? _T_257_89_2 : _GEN_1382;
  wire  _GEN_1387 = 8'h59 == io_fetchQuery_index ? _T_257_89_3 : _GEN_1383;
  wire  _GEN_1388 = 8'h5a == io_fetchQuery_index ? _T_257_90_0 : _GEN_1384;
  wire  _GEN_1389 = 8'h5a == io_fetchQuery_index ? _T_257_90_1 : _GEN_1385;
  wire  _GEN_1390 = 8'h5a == io_fetchQuery_index ? _T_257_90_2 : _GEN_1386;
  wire  _GEN_1391 = 8'h5a == io_fetchQuery_index ? _T_257_90_3 : _GEN_1387;
  wire  _GEN_1392 = 8'h5b == io_fetchQuery_index ? _T_257_91_0 : _GEN_1388;
  wire  _GEN_1393 = 8'h5b == io_fetchQuery_index ? _T_257_91_1 : _GEN_1389;
  wire  _GEN_1394 = 8'h5b == io_fetchQuery_index ? _T_257_91_2 : _GEN_1390;
  wire  _GEN_1395 = 8'h5b == io_fetchQuery_index ? _T_257_91_3 : _GEN_1391;
  wire  _GEN_1396 = 8'h5c == io_fetchQuery_index ? _T_257_92_0 : _GEN_1392;
  wire  _GEN_1397 = 8'h5c == io_fetchQuery_index ? _T_257_92_1 : _GEN_1393;
  wire  _GEN_1398 = 8'h5c == io_fetchQuery_index ? _T_257_92_2 : _GEN_1394;
  wire  _GEN_1399 = 8'h5c == io_fetchQuery_index ? _T_257_92_3 : _GEN_1395;
  wire  _GEN_1400 = 8'h5d == io_fetchQuery_index ? _T_257_93_0 : _GEN_1396;
  wire  _GEN_1401 = 8'h5d == io_fetchQuery_index ? _T_257_93_1 : _GEN_1397;
  wire  _GEN_1402 = 8'h5d == io_fetchQuery_index ? _T_257_93_2 : _GEN_1398;
  wire  _GEN_1403 = 8'h5d == io_fetchQuery_index ? _T_257_93_3 : _GEN_1399;
  wire  _GEN_1404 = 8'h5e == io_fetchQuery_index ? _T_257_94_0 : _GEN_1400;
  wire  _GEN_1405 = 8'h5e == io_fetchQuery_index ? _T_257_94_1 : _GEN_1401;
  wire  _GEN_1406 = 8'h5e == io_fetchQuery_index ? _T_257_94_2 : _GEN_1402;
  wire  _GEN_1407 = 8'h5e == io_fetchQuery_index ? _T_257_94_3 : _GEN_1403;
  wire  _GEN_1408 = 8'h5f == io_fetchQuery_index ? _T_257_95_0 : _GEN_1404;
  wire  _GEN_1409 = 8'h5f == io_fetchQuery_index ? _T_257_95_1 : _GEN_1405;
  wire  _GEN_1410 = 8'h5f == io_fetchQuery_index ? _T_257_95_2 : _GEN_1406;
  wire  _GEN_1411 = 8'h5f == io_fetchQuery_index ? _T_257_95_3 : _GEN_1407;
  wire  _GEN_1412 = 8'h60 == io_fetchQuery_index ? _T_257_96_0 : _GEN_1408;
  wire  _GEN_1413 = 8'h60 == io_fetchQuery_index ? _T_257_96_1 : _GEN_1409;
  wire  _GEN_1414 = 8'h60 == io_fetchQuery_index ? _T_257_96_2 : _GEN_1410;
  wire  _GEN_1415 = 8'h60 == io_fetchQuery_index ? _T_257_96_3 : _GEN_1411;
  wire  _GEN_1416 = 8'h61 == io_fetchQuery_index ? _T_257_97_0 : _GEN_1412;
  wire  _GEN_1417 = 8'h61 == io_fetchQuery_index ? _T_257_97_1 : _GEN_1413;
  wire  _GEN_1418 = 8'h61 == io_fetchQuery_index ? _T_257_97_2 : _GEN_1414;
  wire  _GEN_1419 = 8'h61 == io_fetchQuery_index ? _T_257_97_3 : _GEN_1415;
  wire  _GEN_1420 = 8'h62 == io_fetchQuery_index ? _T_257_98_0 : _GEN_1416;
  wire  _GEN_1421 = 8'h62 == io_fetchQuery_index ? _T_257_98_1 : _GEN_1417;
  wire  _GEN_1422 = 8'h62 == io_fetchQuery_index ? _T_257_98_2 : _GEN_1418;
  wire  _GEN_1423 = 8'h62 == io_fetchQuery_index ? _T_257_98_3 : _GEN_1419;
  wire  _GEN_1424 = 8'h63 == io_fetchQuery_index ? _T_257_99_0 : _GEN_1420;
  wire  _GEN_1425 = 8'h63 == io_fetchQuery_index ? _T_257_99_1 : _GEN_1421;
  wire  _GEN_1426 = 8'h63 == io_fetchQuery_index ? _T_257_99_2 : _GEN_1422;
  wire  _GEN_1427 = 8'h63 == io_fetchQuery_index ? _T_257_99_3 : _GEN_1423;
  wire  _GEN_1428 = 8'h64 == io_fetchQuery_index ? _T_257_100_0 : _GEN_1424;
  wire  _GEN_1429 = 8'h64 == io_fetchQuery_index ? _T_257_100_1 : _GEN_1425;
  wire  _GEN_1430 = 8'h64 == io_fetchQuery_index ? _T_257_100_2 : _GEN_1426;
  wire  _GEN_1431 = 8'h64 == io_fetchQuery_index ? _T_257_100_3 : _GEN_1427;
  wire  _GEN_1432 = 8'h65 == io_fetchQuery_index ? _T_257_101_0 : _GEN_1428;
  wire  _GEN_1433 = 8'h65 == io_fetchQuery_index ? _T_257_101_1 : _GEN_1429;
  wire  _GEN_1434 = 8'h65 == io_fetchQuery_index ? _T_257_101_2 : _GEN_1430;
  wire  _GEN_1435 = 8'h65 == io_fetchQuery_index ? _T_257_101_3 : _GEN_1431;
  wire  _GEN_1436 = 8'h66 == io_fetchQuery_index ? _T_257_102_0 : _GEN_1432;
  wire  _GEN_1437 = 8'h66 == io_fetchQuery_index ? _T_257_102_1 : _GEN_1433;
  wire  _GEN_1438 = 8'h66 == io_fetchQuery_index ? _T_257_102_2 : _GEN_1434;
  wire  _GEN_1439 = 8'h66 == io_fetchQuery_index ? _T_257_102_3 : _GEN_1435;
  wire  _GEN_1440 = 8'h67 == io_fetchQuery_index ? _T_257_103_0 : _GEN_1436;
  wire  _GEN_1441 = 8'h67 == io_fetchQuery_index ? _T_257_103_1 : _GEN_1437;
  wire  _GEN_1442 = 8'h67 == io_fetchQuery_index ? _T_257_103_2 : _GEN_1438;
  wire  _GEN_1443 = 8'h67 == io_fetchQuery_index ? _T_257_103_3 : _GEN_1439;
  wire  _GEN_1444 = 8'h68 == io_fetchQuery_index ? _T_257_104_0 : _GEN_1440;
  wire  _GEN_1445 = 8'h68 == io_fetchQuery_index ? _T_257_104_1 : _GEN_1441;
  wire  _GEN_1446 = 8'h68 == io_fetchQuery_index ? _T_257_104_2 : _GEN_1442;
  wire  _GEN_1447 = 8'h68 == io_fetchQuery_index ? _T_257_104_3 : _GEN_1443;
  wire  _GEN_1448 = 8'h69 == io_fetchQuery_index ? _T_257_105_0 : _GEN_1444;
  wire  _GEN_1449 = 8'h69 == io_fetchQuery_index ? _T_257_105_1 : _GEN_1445;
  wire  _GEN_1450 = 8'h69 == io_fetchQuery_index ? _T_257_105_2 : _GEN_1446;
  wire  _GEN_1451 = 8'h69 == io_fetchQuery_index ? _T_257_105_3 : _GEN_1447;
  wire  _GEN_1452 = 8'h6a == io_fetchQuery_index ? _T_257_106_0 : _GEN_1448;
  wire  _GEN_1453 = 8'h6a == io_fetchQuery_index ? _T_257_106_1 : _GEN_1449;
  wire  _GEN_1454 = 8'h6a == io_fetchQuery_index ? _T_257_106_2 : _GEN_1450;
  wire  _GEN_1455 = 8'h6a == io_fetchQuery_index ? _T_257_106_3 : _GEN_1451;
  wire  _GEN_1456 = 8'h6b == io_fetchQuery_index ? _T_257_107_0 : _GEN_1452;
  wire  _GEN_1457 = 8'h6b == io_fetchQuery_index ? _T_257_107_1 : _GEN_1453;
  wire  _GEN_1458 = 8'h6b == io_fetchQuery_index ? _T_257_107_2 : _GEN_1454;
  wire  _GEN_1459 = 8'h6b == io_fetchQuery_index ? _T_257_107_3 : _GEN_1455;
  wire  _GEN_1460 = 8'h6c == io_fetchQuery_index ? _T_257_108_0 : _GEN_1456;
  wire  _GEN_1461 = 8'h6c == io_fetchQuery_index ? _T_257_108_1 : _GEN_1457;
  wire  _GEN_1462 = 8'h6c == io_fetchQuery_index ? _T_257_108_2 : _GEN_1458;
  wire  _GEN_1463 = 8'h6c == io_fetchQuery_index ? _T_257_108_3 : _GEN_1459;
  wire  _GEN_1464 = 8'h6d == io_fetchQuery_index ? _T_257_109_0 : _GEN_1460;
  wire  _GEN_1465 = 8'h6d == io_fetchQuery_index ? _T_257_109_1 : _GEN_1461;
  wire  _GEN_1466 = 8'h6d == io_fetchQuery_index ? _T_257_109_2 : _GEN_1462;
  wire  _GEN_1467 = 8'h6d == io_fetchQuery_index ? _T_257_109_3 : _GEN_1463;
  wire  _GEN_1468 = 8'h6e == io_fetchQuery_index ? _T_257_110_0 : _GEN_1464;
  wire  _GEN_1469 = 8'h6e == io_fetchQuery_index ? _T_257_110_1 : _GEN_1465;
  wire  _GEN_1470 = 8'h6e == io_fetchQuery_index ? _T_257_110_2 : _GEN_1466;
  wire  _GEN_1471 = 8'h6e == io_fetchQuery_index ? _T_257_110_3 : _GEN_1467;
  wire  _GEN_1472 = 8'h6f == io_fetchQuery_index ? _T_257_111_0 : _GEN_1468;
  wire  _GEN_1473 = 8'h6f == io_fetchQuery_index ? _T_257_111_1 : _GEN_1469;
  wire  _GEN_1474 = 8'h6f == io_fetchQuery_index ? _T_257_111_2 : _GEN_1470;
  wire  _GEN_1475 = 8'h6f == io_fetchQuery_index ? _T_257_111_3 : _GEN_1471;
  wire  _GEN_1476 = 8'h70 == io_fetchQuery_index ? _T_257_112_0 : _GEN_1472;
  wire  _GEN_1477 = 8'h70 == io_fetchQuery_index ? _T_257_112_1 : _GEN_1473;
  wire  _GEN_1478 = 8'h70 == io_fetchQuery_index ? _T_257_112_2 : _GEN_1474;
  wire  _GEN_1479 = 8'h70 == io_fetchQuery_index ? _T_257_112_3 : _GEN_1475;
  wire  _GEN_1480 = 8'h71 == io_fetchQuery_index ? _T_257_113_0 : _GEN_1476;
  wire  _GEN_1481 = 8'h71 == io_fetchQuery_index ? _T_257_113_1 : _GEN_1477;
  wire  _GEN_1482 = 8'h71 == io_fetchQuery_index ? _T_257_113_2 : _GEN_1478;
  wire  _GEN_1483 = 8'h71 == io_fetchQuery_index ? _T_257_113_3 : _GEN_1479;
  wire  _GEN_1484 = 8'h72 == io_fetchQuery_index ? _T_257_114_0 : _GEN_1480;
  wire  _GEN_1485 = 8'h72 == io_fetchQuery_index ? _T_257_114_1 : _GEN_1481;
  wire  _GEN_1486 = 8'h72 == io_fetchQuery_index ? _T_257_114_2 : _GEN_1482;
  wire  _GEN_1487 = 8'h72 == io_fetchQuery_index ? _T_257_114_3 : _GEN_1483;
  wire  _GEN_1488 = 8'h73 == io_fetchQuery_index ? _T_257_115_0 : _GEN_1484;
  wire  _GEN_1489 = 8'h73 == io_fetchQuery_index ? _T_257_115_1 : _GEN_1485;
  wire  _GEN_1490 = 8'h73 == io_fetchQuery_index ? _T_257_115_2 : _GEN_1486;
  wire  _GEN_1491 = 8'h73 == io_fetchQuery_index ? _T_257_115_3 : _GEN_1487;
  wire  _GEN_1492 = 8'h74 == io_fetchQuery_index ? _T_257_116_0 : _GEN_1488;
  wire  _GEN_1493 = 8'h74 == io_fetchQuery_index ? _T_257_116_1 : _GEN_1489;
  wire  _GEN_1494 = 8'h74 == io_fetchQuery_index ? _T_257_116_2 : _GEN_1490;
  wire  _GEN_1495 = 8'h74 == io_fetchQuery_index ? _T_257_116_3 : _GEN_1491;
  wire  _GEN_1496 = 8'h75 == io_fetchQuery_index ? _T_257_117_0 : _GEN_1492;
  wire  _GEN_1497 = 8'h75 == io_fetchQuery_index ? _T_257_117_1 : _GEN_1493;
  wire  _GEN_1498 = 8'h75 == io_fetchQuery_index ? _T_257_117_2 : _GEN_1494;
  wire  _GEN_1499 = 8'h75 == io_fetchQuery_index ? _T_257_117_3 : _GEN_1495;
  wire  _GEN_1500 = 8'h76 == io_fetchQuery_index ? _T_257_118_0 : _GEN_1496;
  wire  _GEN_1501 = 8'h76 == io_fetchQuery_index ? _T_257_118_1 : _GEN_1497;
  wire  _GEN_1502 = 8'h76 == io_fetchQuery_index ? _T_257_118_2 : _GEN_1498;
  wire  _GEN_1503 = 8'h76 == io_fetchQuery_index ? _T_257_118_3 : _GEN_1499;
  wire  _GEN_1504 = 8'h77 == io_fetchQuery_index ? _T_257_119_0 : _GEN_1500;
  wire  _GEN_1505 = 8'h77 == io_fetchQuery_index ? _T_257_119_1 : _GEN_1501;
  wire  _GEN_1506 = 8'h77 == io_fetchQuery_index ? _T_257_119_2 : _GEN_1502;
  wire  _GEN_1507 = 8'h77 == io_fetchQuery_index ? _T_257_119_3 : _GEN_1503;
  wire  _GEN_1508 = 8'h78 == io_fetchQuery_index ? _T_257_120_0 : _GEN_1504;
  wire  _GEN_1509 = 8'h78 == io_fetchQuery_index ? _T_257_120_1 : _GEN_1505;
  wire  _GEN_1510 = 8'h78 == io_fetchQuery_index ? _T_257_120_2 : _GEN_1506;
  wire  _GEN_1511 = 8'h78 == io_fetchQuery_index ? _T_257_120_3 : _GEN_1507;
  wire  _GEN_1512 = 8'h79 == io_fetchQuery_index ? _T_257_121_0 : _GEN_1508;
  wire  _GEN_1513 = 8'h79 == io_fetchQuery_index ? _T_257_121_1 : _GEN_1509;
  wire  _GEN_1514 = 8'h79 == io_fetchQuery_index ? _T_257_121_2 : _GEN_1510;
  wire  _GEN_1515 = 8'h79 == io_fetchQuery_index ? _T_257_121_3 : _GEN_1511;
  wire  _GEN_1516 = 8'h7a == io_fetchQuery_index ? _T_257_122_0 : _GEN_1512;
  wire  _GEN_1517 = 8'h7a == io_fetchQuery_index ? _T_257_122_1 : _GEN_1513;
  wire  _GEN_1518 = 8'h7a == io_fetchQuery_index ? _T_257_122_2 : _GEN_1514;
  wire  _GEN_1519 = 8'h7a == io_fetchQuery_index ? _T_257_122_3 : _GEN_1515;
  wire  _GEN_1520 = 8'h7b == io_fetchQuery_index ? _T_257_123_0 : _GEN_1516;
  wire  _GEN_1521 = 8'h7b == io_fetchQuery_index ? _T_257_123_1 : _GEN_1517;
  wire  _GEN_1522 = 8'h7b == io_fetchQuery_index ? _T_257_123_2 : _GEN_1518;
  wire  _GEN_1523 = 8'h7b == io_fetchQuery_index ? _T_257_123_3 : _GEN_1519;
  wire  _GEN_1524 = 8'h7c == io_fetchQuery_index ? _T_257_124_0 : _GEN_1520;
  wire  _GEN_1525 = 8'h7c == io_fetchQuery_index ? _T_257_124_1 : _GEN_1521;
  wire  _GEN_1526 = 8'h7c == io_fetchQuery_index ? _T_257_124_2 : _GEN_1522;
  wire  _GEN_1527 = 8'h7c == io_fetchQuery_index ? _T_257_124_3 : _GEN_1523;
  wire  _GEN_1528 = 8'h7d == io_fetchQuery_index ? _T_257_125_0 : _GEN_1524;
  wire  _GEN_1529 = 8'h7d == io_fetchQuery_index ? _T_257_125_1 : _GEN_1525;
  wire  _GEN_1530 = 8'h7d == io_fetchQuery_index ? _T_257_125_2 : _GEN_1526;
  wire  _GEN_1531 = 8'h7d == io_fetchQuery_index ? _T_257_125_3 : _GEN_1527;
  wire  _GEN_1532 = 8'h7e == io_fetchQuery_index ? _T_257_126_0 : _GEN_1528;
  wire  _GEN_1533 = 8'h7e == io_fetchQuery_index ? _T_257_126_1 : _GEN_1529;
  wire  _GEN_1534 = 8'h7e == io_fetchQuery_index ? _T_257_126_2 : _GEN_1530;
  wire  _GEN_1535 = 8'h7e == io_fetchQuery_index ? _T_257_126_3 : _GEN_1531;
  wire  _GEN_1536 = 8'h7f == io_fetchQuery_index ? _T_257_127_0 : _GEN_1532;
  wire  _GEN_1537 = 8'h7f == io_fetchQuery_index ? _T_257_127_1 : _GEN_1533;
  wire  _GEN_1538 = 8'h7f == io_fetchQuery_index ? _T_257_127_2 : _GEN_1534;
  wire  _GEN_1539 = 8'h7f == io_fetchQuery_index ? _T_257_127_3 : _GEN_1535;
  wire  _GEN_1540 = 8'h80 == io_fetchQuery_index ? _T_257_128_0 : _GEN_1536;
  wire  _GEN_1541 = 8'h80 == io_fetchQuery_index ? _T_257_128_1 : _GEN_1537;
  wire  _GEN_1542 = 8'h80 == io_fetchQuery_index ? _T_257_128_2 : _GEN_1538;
  wire  _GEN_1543 = 8'h80 == io_fetchQuery_index ? _T_257_128_3 : _GEN_1539;
  wire  _GEN_1544 = 8'h81 == io_fetchQuery_index ? _T_257_129_0 : _GEN_1540;
  wire  _GEN_1545 = 8'h81 == io_fetchQuery_index ? _T_257_129_1 : _GEN_1541;
  wire  _GEN_1546 = 8'h81 == io_fetchQuery_index ? _T_257_129_2 : _GEN_1542;
  wire  _GEN_1547 = 8'h81 == io_fetchQuery_index ? _T_257_129_3 : _GEN_1543;
  wire  _GEN_1548 = 8'h82 == io_fetchQuery_index ? _T_257_130_0 : _GEN_1544;
  wire  _GEN_1549 = 8'h82 == io_fetchQuery_index ? _T_257_130_1 : _GEN_1545;
  wire  _GEN_1550 = 8'h82 == io_fetchQuery_index ? _T_257_130_2 : _GEN_1546;
  wire  _GEN_1551 = 8'h82 == io_fetchQuery_index ? _T_257_130_3 : _GEN_1547;
  wire  _GEN_1552 = 8'h83 == io_fetchQuery_index ? _T_257_131_0 : _GEN_1548;
  wire  _GEN_1553 = 8'h83 == io_fetchQuery_index ? _T_257_131_1 : _GEN_1549;
  wire  _GEN_1554 = 8'h83 == io_fetchQuery_index ? _T_257_131_2 : _GEN_1550;
  wire  _GEN_1555 = 8'h83 == io_fetchQuery_index ? _T_257_131_3 : _GEN_1551;
  wire  _GEN_1556 = 8'h84 == io_fetchQuery_index ? _T_257_132_0 : _GEN_1552;
  wire  _GEN_1557 = 8'h84 == io_fetchQuery_index ? _T_257_132_1 : _GEN_1553;
  wire  _GEN_1558 = 8'h84 == io_fetchQuery_index ? _T_257_132_2 : _GEN_1554;
  wire  _GEN_1559 = 8'h84 == io_fetchQuery_index ? _T_257_132_3 : _GEN_1555;
  wire  _GEN_1560 = 8'h85 == io_fetchQuery_index ? _T_257_133_0 : _GEN_1556;
  wire  _GEN_1561 = 8'h85 == io_fetchQuery_index ? _T_257_133_1 : _GEN_1557;
  wire  _GEN_1562 = 8'h85 == io_fetchQuery_index ? _T_257_133_2 : _GEN_1558;
  wire  _GEN_1563 = 8'h85 == io_fetchQuery_index ? _T_257_133_3 : _GEN_1559;
  wire  _GEN_1564 = 8'h86 == io_fetchQuery_index ? _T_257_134_0 : _GEN_1560;
  wire  _GEN_1565 = 8'h86 == io_fetchQuery_index ? _T_257_134_1 : _GEN_1561;
  wire  _GEN_1566 = 8'h86 == io_fetchQuery_index ? _T_257_134_2 : _GEN_1562;
  wire  _GEN_1567 = 8'h86 == io_fetchQuery_index ? _T_257_134_3 : _GEN_1563;
  wire  _GEN_1568 = 8'h87 == io_fetchQuery_index ? _T_257_135_0 : _GEN_1564;
  wire  _GEN_1569 = 8'h87 == io_fetchQuery_index ? _T_257_135_1 : _GEN_1565;
  wire  _GEN_1570 = 8'h87 == io_fetchQuery_index ? _T_257_135_2 : _GEN_1566;
  wire  _GEN_1571 = 8'h87 == io_fetchQuery_index ? _T_257_135_3 : _GEN_1567;
  wire  _GEN_1572 = 8'h88 == io_fetchQuery_index ? _T_257_136_0 : _GEN_1568;
  wire  _GEN_1573 = 8'h88 == io_fetchQuery_index ? _T_257_136_1 : _GEN_1569;
  wire  _GEN_1574 = 8'h88 == io_fetchQuery_index ? _T_257_136_2 : _GEN_1570;
  wire  _GEN_1575 = 8'h88 == io_fetchQuery_index ? _T_257_136_3 : _GEN_1571;
  wire  _GEN_1576 = 8'h89 == io_fetchQuery_index ? _T_257_137_0 : _GEN_1572;
  wire  _GEN_1577 = 8'h89 == io_fetchQuery_index ? _T_257_137_1 : _GEN_1573;
  wire  _GEN_1578 = 8'h89 == io_fetchQuery_index ? _T_257_137_2 : _GEN_1574;
  wire  _GEN_1579 = 8'h89 == io_fetchQuery_index ? _T_257_137_3 : _GEN_1575;
  wire  _GEN_1580 = 8'h8a == io_fetchQuery_index ? _T_257_138_0 : _GEN_1576;
  wire  _GEN_1581 = 8'h8a == io_fetchQuery_index ? _T_257_138_1 : _GEN_1577;
  wire  _GEN_1582 = 8'h8a == io_fetchQuery_index ? _T_257_138_2 : _GEN_1578;
  wire  _GEN_1583 = 8'h8a == io_fetchQuery_index ? _T_257_138_3 : _GEN_1579;
  wire  _GEN_1584 = 8'h8b == io_fetchQuery_index ? _T_257_139_0 : _GEN_1580;
  wire  _GEN_1585 = 8'h8b == io_fetchQuery_index ? _T_257_139_1 : _GEN_1581;
  wire  _GEN_1586 = 8'h8b == io_fetchQuery_index ? _T_257_139_2 : _GEN_1582;
  wire  _GEN_1587 = 8'h8b == io_fetchQuery_index ? _T_257_139_3 : _GEN_1583;
  wire  _GEN_1588 = 8'h8c == io_fetchQuery_index ? _T_257_140_0 : _GEN_1584;
  wire  _GEN_1589 = 8'h8c == io_fetchQuery_index ? _T_257_140_1 : _GEN_1585;
  wire  _GEN_1590 = 8'h8c == io_fetchQuery_index ? _T_257_140_2 : _GEN_1586;
  wire  _GEN_1591 = 8'h8c == io_fetchQuery_index ? _T_257_140_3 : _GEN_1587;
  wire  _GEN_1592 = 8'h8d == io_fetchQuery_index ? _T_257_141_0 : _GEN_1588;
  wire  _GEN_1593 = 8'h8d == io_fetchQuery_index ? _T_257_141_1 : _GEN_1589;
  wire  _GEN_1594 = 8'h8d == io_fetchQuery_index ? _T_257_141_2 : _GEN_1590;
  wire  _GEN_1595 = 8'h8d == io_fetchQuery_index ? _T_257_141_3 : _GEN_1591;
  wire  _GEN_1596 = 8'h8e == io_fetchQuery_index ? _T_257_142_0 : _GEN_1592;
  wire  _GEN_1597 = 8'h8e == io_fetchQuery_index ? _T_257_142_1 : _GEN_1593;
  wire  _GEN_1598 = 8'h8e == io_fetchQuery_index ? _T_257_142_2 : _GEN_1594;
  wire  _GEN_1599 = 8'h8e == io_fetchQuery_index ? _T_257_142_3 : _GEN_1595;
  wire  _GEN_1600 = 8'h8f == io_fetchQuery_index ? _T_257_143_0 : _GEN_1596;
  wire  _GEN_1601 = 8'h8f == io_fetchQuery_index ? _T_257_143_1 : _GEN_1597;
  wire  _GEN_1602 = 8'h8f == io_fetchQuery_index ? _T_257_143_2 : _GEN_1598;
  wire  _GEN_1603 = 8'h8f == io_fetchQuery_index ? _T_257_143_3 : _GEN_1599;
  wire  _GEN_1604 = 8'h90 == io_fetchQuery_index ? _T_257_144_0 : _GEN_1600;
  wire  _GEN_1605 = 8'h90 == io_fetchQuery_index ? _T_257_144_1 : _GEN_1601;
  wire  _GEN_1606 = 8'h90 == io_fetchQuery_index ? _T_257_144_2 : _GEN_1602;
  wire  _GEN_1607 = 8'h90 == io_fetchQuery_index ? _T_257_144_3 : _GEN_1603;
  wire  _GEN_1608 = 8'h91 == io_fetchQuery_index ? _T_257_145_0 : _GEN_1604;
  wire  _GEN_1609 = 8'h91 == io_fetchQuery_index ? _T_257_145_1 : _GEN_1605;
  wire  _GEN_1610 = 8'h91 == io_fetchQuery_index ? _T_257_145_2 : _GEN_1606;
  wire  _GEN_1611 = 8'h91 == io_fetchQuery_index ? _T_257_145_3 : _GEN_1607;
  wire  _GEN_1612 = 8'h92 == io_fetchQuery_index ? _T_257_146_0 : _GEN_1608;
  wire  _GEN_1613 = 8'h92 == io_fetchQuery_index ? _T_257_146_1 : _GEN_1609;
  wire  _GEN_1614 = 8'h92 == io_fetchQuery_index ? _T_257_146_2 : _GEN_1610;
  wire  _GEN_1615 = 8'h92 == io_fetchQuery_index ? _T_257_146_3 : _GEN_1611;
  wire  _GEN_1616 = 8'h93 == io_fetchQuery_index ? _T_257_147_0 : _GEN_1612;
  wire  _GEN_1617 = 8'h93 == io_fetchQuery_index ? _T_257_147_1 : _GEN_1613;
  wire  _GEN_1618 = 8'h93 == io_fetchQuery_index ? _T_257_147_2 : _GEN_1614;
  wire  _GEN_1619 = 8'h93 == io_fetchQuery_index ? _T_257_147_3 : _GEN_1615;
  wire  _GEN_1620 = 8'h94 == io_fetchQuery_index ? _T_257_148_0 : _GEN_1616;
  wire  _GEN_1621 = 8'h94 == io_fetchQuery_index ? _T_257_148_1 : _GEN_1617;
  wire  _GEN_1622 = 8'h94 == io_fetchQuery_index ? _T_257_148_2 : _GEN_1618;
  wire  _GEN_1623 = 8'h94 == io_fetchQuery_index ? _T_257_148_3 : _GEN_1619;
  wire  _GEN_1624 = 8'h95 == io_fetchQuery_index ? _T_257_149_0 : _GEN_1620;
  wire  _GEN_1625 = 8'h95 == io_fetchQuery_index ? _T_257_149_1 : _GEN_1621;
  wire  _GEN_1626 = 8'h95 == io_fetchQuery_index ? _T_257_149_2 : _GEN_1622;
  wire  _GEN_1627 = 8'h95 == io_fetchQuery_index ? _T_257_149_3 : _GEN_1623;
  wire  _GEN_1628 = 8'h96 == io_fetchQuery_index ? _T_257_150_0 : _GEN_1624;
  wire  _GEN_1629 = 8'h96 == io_fetchQuery_index ? _T_257_150_1 : _GEN_1625;
  wire  _GEN_1630 = 8'h96 == io_fetchQuery_index ? _T_257_150_2 : _GEN_1626;
  wire  _GEN_1631 = 8'h96 == io_fetchQuery_index ? _T_257_150_3 : _GEN_1627;
  wire  _GEN_1632 = 8'h97 == io_fetchQuery_index ? _T_257_151_0 : _GEN_1628;
  wire  _GEN_1633 = 8'h97 == io_fetchQuery_index ? _T_257_151_1 : _GEN_1629;
  wire  _GEN_1634 = 8'h97 == io_fetchQuery_index ? _T_257_151_2 : _GEN_1630;
  wire  _GEN_1635 = 8'h97 == io_fetchQuery_index ? _T_257_151_3 : _GEN_1631;
  wire  _GEN_1636 = 8'h98 == io_fetchQuery_index ? _T_257_152_0 : _GEN_1632;
  wire  _GEN_1637 = 8'h98 == io_fetchQuery_index ? _T_257_152_1 : _GEN_1633;
  wire  _GEN_1638 = 8'h98 == io_fetchQuery_index ? _T_257_152_2 : _GEN_1634;
  wire  _GEN_1639 = 8'h98 == io_fetchQuery_index ? _T_257_152_3 : _GEN_1635;
  wire  _GEN_1640 = 8'h99 == io_fetchQuery_index ? _T_257_153_0 : _GEN_1636;
  wire  _GEN_1641 = 8'h99 == io_fetchQuery_index ? _T_257_153_1 : _GEN_1637;
  wire  _GEN_1642 = 8'h99 == io_fetchQuery_index ? _T_257_153_2 : _GEN_1638;
  wire  _GEN_1643 = 8'h99 == io_fetchQuery_index ? _T_257_153_3 : _GEN_1639;
  wire  _GEN_1644 = 8'h9a == io_fetchQuery_index ? _T_257_154_0 : _GEN_1640;
  wire  _GEN_1645 = 8'h9a == io_fetchQuery_index ? _T_257_154_1 : _GEN_1641;
  wire  _GEN_1646 = 8'h9a == io_fetchQuery_index ? _T_257_154_2 : _GEN_1642;
  wire  _GEN_1647 = 8'h9a == io_fetchQuery_index ? _T_257_154_3 : _GEN_1643;
  wire  _GEN_1648 = 8'h9b == io_fetchQuery_index ? _T_257_155_0 : _GEN_1644;
  wire  _GEN_1649 = 8'h9b == io_fetchQuery_index ? _T_257_155_1 : _GEN_1645;
  wire  _GEN_1650 = 8'h9b == io_fetchQuery_index ? _T_257_155_2 : _GEN_1646;
  wire  _GEN_1651 = 8'h9b == io_fetchQuery_index ? _T_257_155_3 : _GEN_1647;
  wire  _GEN_1652 = 8'h9c == io_fetchQuery_index ? _T_257_156_0 : _GEN_1648;
  wire  _GEN_1653 = 8'h9c == io_fetchQuery_index ? _T_257_156_1 : _GEN_1649;
  wire  _GEN_1654 = 8'h9c == io_fetchQuery_index ? _T_257_156_2 : _GEN_1650;
  wire  _GEN_1655 = 8'h9c == io_fetchQuery_index ? _T_257_156_3 : _GEN_1651;
  wire  _GEN_1656 = 8'h9d == io_fetchQuery_index ? _T_257_157_0 : _GEN_1652;
  wire  _GEN_1657 = 8'h9d == io_fetchQuery_index ? _T_257_157_1 : _GEN_1653;
  wire  _GEN_1658 = 8'h9d == io_fetchQuery_index ? _T_257_157_2 : _GEN_1654;
  wire  _GEN_1659 = 8'h9d == io_fetchQuery_index ? _T_257_157_3 : _GEN_1655;
  wire  _GEN_1660 = 8'h9e == io_fetchQuery_index ? _T_257_158_0 : _GEN_1656;
  wire  _GEN_1661 = 8'h9e == io_fetchQuery_index ? _T_257_158_1 : _GEN_1657;
  wire  _GEN_1662 = 8'h9e == io_fetchQuery_index ? _T_257_158_2 : _GEN_1658;
  wire  _GEN_1663 = 8'h9e == io_fetchQuery_index ? _T_257_158_3 : _GEN_1659;
  wire  _GEN_1664 = 8'h9f == io_fetchQuery_index ? _T_257_159_0 : _GEN_1660;
  wire  _GEN_1665 = 8'h9f == io_fetchQuery_index ? _T_257_159_1 : _GEN_1661;
  wire  _GEN_1666 = 8'h9f == io_fetchQuery_index ? _T_257_159_2 : _GEN_1662;
  wire  _GEN_1667 = 8'h9f == io_fetchQuery_index ? _T_257_159_3 : _GEN_1663;
  wire  _GEN_1668 = 8'ha0 == io_fetchQuery_index ? _T_257_160_0 : _GEN_1664;
  wire  _GEN_1669 = 8'ha0 == io_fetchQuery_index ? _T_257_160_1 : _GEN_1665;
  wire  _GEN_1670 = 8'ha0 == io_fetchQuery_index ? _T_257_160_2 : _GEN_1666;
  wire  _GEN_1671 = 8'ha0 == io_fetchQuery_index ? _T_257_160_3 : _GEN_1667;
  wire  _GEN_1672 = 8'ha1 == io_fetchQuery_index ? _T_257_161_0 : _GEN_1668;
  wire  _GEN_1673 = 8'ha1 == io_fetchQuery_index ? _T_257_161_1 : _GEN_1669;
  wire  _GEN_1674 = 8'ha1 == io_fetchQuery_index ? _T_257_161_2 : _GEN_1670;
  wire  _GEN_1675 = 8'ha1 == io_fetchQuery_index ? _T_257_161_3 : _GEN_1671;
  wire  _GEN_1676 = 8'ha2 == io_fetchQuery_index ? _T_257_162_0 : _GEN_1672;
  wire  _GEN_1677 = 8'ha2 == io_fetchQuery_index ? _T_257_162_1 : _GEN_1673;
  wire  _GEN_1678 = 8'ha2 == io_fetchQuery_index ? _T_257_162_2 : _GEN_1674;
  wire  _GEN_1679 = 8'ha2 == io_fetchQuery_index ? _T_257_162_3 : _GEN_1675;
  wire  _GEN_1680 = 8'ha3 == io_fetchQuery_index ? _T_257_163_0 : _GEN_1676;
  wire  _GEN_1681 = 8'ha3 == io_fetchQuery_index ? _T_257_163_1 : _GEN_1677;
  wire  _GEN_1682 = 8'ha3 == io_fetchQuery_index ? _T_257_163_2 : _GEN_1678;
  wire  _GEN_1683 = 8'ha3 == io_fetchQuery_index ? _T_257_163_3 : _GEN_1679;
  wire  _GEN_1684 = 8'ha4 == io_fetchQuery_index ? _T_257_164_0 : _GEN_1680;
  wire  _GEN_1685 = 8'ha4 == io_fetchQuery_index ? _T_257_164_1 : _GEN_1681;
  wire  _GEN_1686 = 8'ha4 == io_fetchQuery_index ? _T_257_164_2 : _GEN_1682;
  wire  _GEN_1687 = 8'ha4 == io_fetchQuery_index ? _T_257_164_3 : _GEN_1683;
  wire  _GEN_1688 = 8'ha5 == io_fetchQuery_index ? _T_257_165_0 : _GEN_1684;
  wire  _GEN_1689 = 8'ha5 == io_fetchQuery_index ? _T_257_165_1 : _GEN_1685;
  wire  _GEN_1690 = 8'ha5 == io_fetchQuery_index ? _T_257_165_2 : _GEN_1686;
  wire  _GEN_1691 = 8'ha5 == io_fetchQuery_index ? _T_257_165_3 : _GEN_1687;
  wire  _GEN_1692 = 8'ha6 == io_fetchQuery_index ? _T_257_166_0 : _GEN_1688;
  wire  _GEN_1693 = 8'ha6 == io_fetchQuery_index ? _T_257_166_1 : _GEN_1689;
  wire  _GEN_1694 = 8'ha6 == io_fetchQuery_index ? _T_257_166_2 : _GEN_1690;
  wire  _GEN_1695 = 8'ha6 == io_fetchQuery_index ? _T_257_166_3 : _GEN_1691;
  wire  _GEN_1696 = 8'ha7 == io_fetchQuery_index ? _T_257_167_0 : _GEN_1692;
  wire  _GEN_1697 = 8'ha7 == io_fetchQuery_index ? _T_257_167_1 : _GEN_1693;
  wire  _GEN_1698 = 8'ha7 == io_fetchQuery_index ? _T_257_167_2 : _GEN_1694;
  wire  _GEN_1699 = 8'ha7 == io_fetchQuery_index ? _T_257_167_3 : _GEN_1695;
  wire  _GEN_1700 = 8'ha8 == io_fetchQuery_index ? _T_257_168_0 : _GEN_1696;
  wire  _GEN_1701 = 8'ha8 == io_fetchQuery_index ? _T_257_168_1 : _GEN_1697;
  wire  _GEN_1702 = 8'ha8 == io_fetchQuery_index ? _T_257_168_2 : _GEN_1698;
  wire  _GEN_1703 = 8'ha8 == io_fetchQuery_index ? _T_257_168_3 : _GEN_1699;
  wire  _GEN_1704 = 8'ha9 == io_fetchQuery_index ? _T_257_169_0 : _GEN_1700;
  wire  _GEN_1705 = 8'ha9 == io_fetchQuery_index ? _T_257_169_1 : _GEN_1701;
  wire  _GEN_1706 = 8'ha9 == io_fetchQuery_index ? _T_257_169_2 : _GEN_1702;
  wire  _GEN_1707 = 8'ha9 == io_fetchQuery_index ? _T_257_169_3 : _GEN_1703;
  wire  _GEN_1708 = 8'haa == io_fetchQuery_index ? _T_257_170_0 : _GEN_1704;
  wire  _GEN_1709 = 8'haa == io_fetchQuery_index ? _T_257_170_1 : _GEN_1705;
  wire  _GEN_1710 = 8'haa == io_fetchQuery_index ? _T_257_170_2 : _GEN_1706;
  wire  _GEN_1711 = 8'haa == io_fetchQuery_index ? _T_257_170_3 : _GEN_1707;
  wire  _GEN_1712 = 8'hab == io_fetchQuery_index ? _T_257_171_0 : _GEN_1708;
  wire  _GEN_1713 = 8'hab == io_fetchQuery_index ? _T_257_171_1 : _GEN_1709;
  wire  _GEN_1714 = 8'hab == io_fetchQuery_index ? _T_257_171_2 : _GEN_1710;
  wire  _GEN_1715 = 8'hab == io_fetchQuery_index ? _T_257_171_3 : _GEN_1711;
  wire  _GEN_1716 = 8'hac == io_fetchQuery_index ? _T_257_172_0 : _GEN_1712;
  wire  _GEN_1717 = 8'hac == io_fetchQuery_index ? _T_257_172_1 : _GEN_1713;
  wire  _GEN_1718 = 8'hac == io_fetchQuery_index ? _T_257_172_2 : _GEN_1714;
  wire  _GEN_1719 = 8'hac == io_fetchQuery_index ? _T_257_172_3 : _GEN_1715;
  wire  _GEN_1720 = 8'had == io_fetchQuery_index ? _T_257_173_0 : _GEN_1716;
  wire  _GEN_1721 = 8'had == io_fetchQuery_index ? _T_257_173_1 : _GEN_1717;
  wire  _GEN_1722 = 8'had == io_fetchQuery_index ? _T_257_173_2 : _GEN_1718;
  wire  _GEN_1723 = 8'had == io_fetchQuery_index ? _T_257_173_3 : _GEN_1719;
  wire  _GEN_1724 = 8'hae == io_fetchQuery_index ? _T_257_174_0 : _GEN_1720;
  wire  _GEN_1725 = 8'hae == io_fetchQuery_index ? _T_257_174_1 : _GEN_1721;
  wire  _GEN_1726 = 8'hae == io_fetchQuery_index ? _T_257_174_2 : _GEN_1722;
  wire  _GEN_1727 = 8'hae == io_fetchQuery_index ? _T_257_174_3 : _GEN_1723;
  wire  _GEN_1728 = 8'haf == io_fetchQuery_index ? _T_257_175_0 : _GEN_1724;
  wire  _GEN_1729 = 8'haf == io_fetchQuery_index ? _T_257_175_1 : _GEN_1725;
  wire  _GEN_1730 = 8'haf == io_fetchQuery_index ? _T_257_175_2 : _GEN_1726;
  wire  _GEN_1731 = 8'haf == io_fetchQuery_index ? _T_257_175_3 : _GEN_1727;
  wire  _GEN_1732 = 8'hb0 == io_fetchQuery_index ? _T_257_176_0 : _GEN_1728;
  wire  _GEN_1733 = 8'hb0 == io_fetchQuery_index ? _T_257_176_1 : _GEN_1729;
  wire  _GEN_1734 = 8'hb0 == io_fetchQuery_index ? _T_257_176_2 : _GEN_1730;
  wire  _GEN_1735 = 8'hb0 == io_fetchQuery_index ? _T_257_176_3 : _GEN_1731;
  wire  _GEN_1736 = 8'hb1 == io_fetchQuery_index ? _T_257_177_0 : _GEN_1732;
  wire  _GEN_1737 = 8'hb1 == io_fetchQuery_index ? _T_257_177_1 : _GEN_1733;
  wire  _GEN_1738 = 8'hb1 == io_fetchQuery_index ? _T_257_177_2 : _GEN_1734;
  wire  _GEN_1739 = 8'hb1 == io_fetchQuery_index ? _T_257_177_3 : _GEN_1735;
  wire  _GEN_1740 = 8'hb2 == io_fetchQuery_index ? _T_257_178_0 : _GEN_1736;
  wire  _GEN_1741 = 8'hb2 == io_fetchQuery_index ? _T_257_178_1 : _GEN_1737;
  wire  _GEN_1742 = 8'hb2 == io_fetchQuery_index ? _T_257_178_2 : _GEN_1738;
  wire  _GEN_1743 = 8'hb2 == io_fetchQuery_index ? _T_257_178_3 : _GEN_1739;
  wire  _GEN_1744 = 8'hb3 == io_fetchQuery_index ? _T_257_179_0 : _GEN_1740;
  wire  _GEN_1745 = 8'hb3 == io_fetchQuery_index ? _T_257_179_1 : _GEN_1741;
  wire  _GEN_1746 = 8'hb3 == io_fetchQuery_index ? _T_257_179_2 : _GEN_1742;
  wire  _GEN_1747 = 8'hb3 == io_fetchQuery_index ? _T_257_179_3 : _GEN_1743;
  wire  _GEN_1748 = 8'hb4 == io_fetchQuery_index ? _T_257_180_0 : _GEN_1744;
  wire  _GEN_1749 = 8'hb4 == io_fetchQuery_index ? _T_257_180_1 : _GEN_1745;
  wire  _GEN_1750 = 8'hb4 == io_fetchQuery_index ? _T_257_180_2 : _GEN_1746;
  wire  _GEN_1751 = 8'hb4 == io_fetchQuery_index ? _T_257_180_3 : _GEN_1747;
  wire  _GEN_1752 = 8'hb5 == io_fetchQuery_index ? _T_257_181_0 : _GEN_1748;
  wire  _GEN_1753 = 8'hb5 == io_fetchQuery_index ? _T_257_181_1 : _GEN_1749;
  wire  _GEN_1754 = 8'hb5 == io_fetchQuery_index ? _T_257_181_2 : _GEN_1750;
  wire  _GEN_1755 = 8'hb5 == io_fetchQuery_index ? _T_257_181_3 : _GEN_1751;
  wire  _GEN_1756 = 8'hb6 == io_fetchQuery_index ? _T_257_182_0 : _GEN_1752;
  wire  _GEN_1757 = 8'hb6 == io_fetchQuery_index ? _T_257_182_1 : _GEN_1753;
  wire  _GEN_1758 = 8'hb6 == io_fetchQuery_index ? _T_257_182_2 : _GEN_1754;
  wire  _GEN_1759 = 8'hb6 == io_fetchQuery_index ? _T_257_182_3 : _GEN_1755;
  wire  _GEN_1760 = 8'hb7 == io_fetchQuery_index ? _T_257_183_0 : _GEN_1756;
  wire  _GEN_1761 = 8'hb7 == io_fetchQuery_index ? _T_257_183_1 : _GEN_1757;
  wire  _GEN_1762 = 8'hb7 == io_fetchQuery_index ? _T_257_183_2 : _GEN_1758;
  wire  _GEN_1763 = 8'hb7 == io_fetchQuery_index ? _T_257_183_3 : _GEN_1759;
  wire  _GEN_1764 = 8'hb8 == io_fetchQuery_index ? _T_257_184_0 : _GEN_1760;
  wire  _GEN_1765 = 8'hb8 == io_fetchQuery_index ? _T_257_184_1 : _GEN_1761;
  wire  _GEN_1766 = 8'hb8 == io_fetchQuery_index ? _T_257_184_2 : _GEN_1762;
  wire  _GEN_1767 = 8'hb8 == io_fetchQuery_index ? _T_257_184_3 : _GEN_1763;
  wire  _GEN_1768 = 8'hb9 == io_fetchQuery_index ? _T_257_185_0 : _GEN_1764;
  wire  _GEN_1769 = 8'hb9 == io_fetchQuery_index ? _T_257_185_1 : _GEN_1765;
  wire  _GEN_1770 = 8'hb9 == io_fetchQuery_index ? _T_257_185_2 : _GEN_1766;
  wire  _GEN_1771 = 8'hb9 == io_fetchQuery_index ? _T_257_185_3 : _GEN_1767;
  wire  _GEN_1772 = 8'hba == io_fetchQuery_index ? _T_257_186_0 : _GEN_1768;
  wire  _GEN_1773 = 8'hba == io_fetchQuery_index ? _T_257_186_1 : _GEN_1769;
  wire  _GEN_1774 = 8'hba == io_fetchQuery_index ? _T_257_186_2 : _GEN_1770;
  wire  _GEN_1775 = 8'hba == io_fetchQuery_index ? _T_257_186_3 : _GEN_1771;
  wire  _GEN_1776 = 8'hbb == io_fetchQuery_index ? _T_257_187_0 : _GEN_1772;
  wire  _GEN_1777 = 8'hbb == io_fetchQuery_index ? _T_257_187_1 : _GEN_1773;
  wire  _GEN_1778 = 8'hbb == io_fetchQuery_index ? _T_257_187_2 : _GEN_1774;
  wire  _GEN_1779 = 8'hbb == io_fetchQuery_index ? _T_257_187_3 : _GEN_1775;
  wire  _GEN_1780 = 8'hbc == io_fetchQuery_index ? _T_257_188_0 : _GEN_1776;
  wire  _GEN_1781 = 8'hbc == io_fetchQuery_index ? _T_257_188_1 : _GEN_1777;
  wire  _GEN_1782 = 8'hbc == io_fetchQuery_index ? _T_257_188_2 : _GEN_1778;
  wire  _GEN_1783 = 8'hbc == io_fetchQuery_index ? _T_257_188_3 : _GEN_1779;
  wire  _GEN_1784 = 8'hbd == io_fetchQuery_index ? _T_257_189_0 : _GEN_1780;
  wire  _GEN_1785 = 8'hbd == io_fetchQuery_index ? _T_257_189_1 : _GEN_1781;
  wire  _GEN_1786 = 8'hbd == io_fetchQuery_index ? _T_257_189_2 : _GEN_1782;
  wire  _GEN_1787 = 8'hbd == io_fetchQuery_index ? _T_257_189_3 : _GEN_1783;
  wire  _GEN_1788 = 8'hbe == io_fetchQuery_index ? _T_257_190_0 : _GEN_1784;
  wire  _GEN_1789 = 8'hbe == io_fetchQuery_index ? _T_257_190_1 : _GEN_1785;
  wire  _GEN_1790 = 8'hbe == io_fetchQuery_index ? _T_257_190_2 : _GEN_1786;
  wire  _GEN_1791 = 8'hbe == io_fetchQuery_index ? _T_257_190_3 : _GEN_1787;
  wire  _GEN_1792 = 8'hbf == io_fetchQuery_index ? _T_257_191_0 : _GEN_1788;
  wire  _GEN_1793 = 8'hbf == io_fetchQuery_index ? _T_257_191_1 : _GEN_1789;
  wire  _GEN_1794 = 8'hbf == io_fetchQuery_index ? _T_257_191_2 : _GEN_1790;
  wire  _GEN_1795 = 8'hbf == io_fetchQuery_index ? _T_257_191_3 : _GEN_1791;
  wire  _GEN_1796 = 8'hc0 == io_fetchQuery_index ? _T_257_192_0 : _GEN_1792;
  wire  _GEN_1797 = 8'hc0 == io_fetchQuery_index ? _T_257_192_1 : _GEN_1793;
  wire  _GEN_1798 = 8'hc0 == io_fetchQuery_index ? _T_257_192_2 : _GEN_1794;
  wire  _GEN_1799 = 8'hc0 == io_fetchQuery_index ? _T_257_192_3 : _GEN_1795;
  wire  _GEN_1800 = 8'hc1 == io_fetchQuery_index ? _T_257_193_0 : _GEN_1796;
  wire  _GEN_1801 = 8'hc1 == io_fetchQuery_index ? _T_257_193_1 : _GEN_1797;
  wire  _GEN_1802 = 8'hc1 == io_fetchQuery_index ? _T_257_193_2 : _GEN_1798;
  wire  _GEN_1803 = 8'hc1 == io_fetchQuery_index ? _T_257_193_3 : _GEN_1799;
  wire  _GEN_1804 = 8'hc2 == io_fetchQuery_index ? _T_257_194_0 : _GEN_1800;
  wire  _GEN_1805 = 8'hc2 == io_fetchQuery_index ? _T_257_194_1 : _GEN_1801;
  wire  _GEN_1806 = 8'hc2 == io_fetchQuery_index ? _T_257_194_2 : _GEN_1802;
  wire  _GEN_1807 = 8'hc2 == io_fetchQuery_index ? _T_257_194_3 : _GEN_1803;
  wire  _GEN_1808 = 8'hc3 == io_fetchQuery_index ? _T_257_195_0 : _GEN_1804;
  wire  _GEN_1809 = 8'hc3 == io_fetchQuery_index ? _T_257_195_1 : _GEN_1805;
  wire  _GEN_1810 = 8'hc3 == io_fetchQuery_index ? _T_257_195_2 : _GEN_1806;
  wire  _GEN_1811 = 8'hc3 == io_fetchQuery_index ? _T_257_195_3 : _GEN_1807;
  wire  _GEN_1812 = 8'hc4 == io_fetchQuery_index ? _T_257_196_0 : _GEN_1808;
  wire  _GEN_1813 = 8'hc4 == io_fetchQuery_index ? _T_257_196_1 : _GEN_1809;
  wire  _GEN_1814 = 8'hc4 == io_fetchQuery_index ? _T_257_196_2 : _GEN_1810;
  wire  _GEN_1815 = 8'hc4 == io_fetchQuery_index ? _T_257_196_3 : _GEN_1811;
  wire  _GEN_1816 = 8'hc5 == io_fetchQuery_index ? _T_257_197_0 : _GEN_1812;
  wire  _GEN_1817 = 8'hc5 == io_fetchQuery_index ? _T_257_197_1 : _GEN_1813;
  wire  _GEN_1818 = 8'hc5 == io_fetchQuery_index ? _T_257_197_2 : _GEN_1814;
  wire  _GEN_1819 = 8'hc5 == io_fetchQuery_index ? _T_257_197_3 : _GEN_1815;
  wire  _GEN_1820 = 8'hc6 == io_fetchQuery_index ? _T_257_198_0 : _GEN_1816;
  wire  _GEN_1821 = 8'hc6 == io_fetchQuery_index ? _T_257_198_1 : _GEN_1817;
  wire  _GEN_1822 = 8'hc6 == io_fetchQuery_index ? _T_257_198_2 : _GEN_1818;
  wire  _GEN_1823 = 8'hc6 == io_fetchQuery_index ? _T_257_198_3 : _GEN_1819;
  wire  _GEN_1824 = 8'hc7 == io_fetchQuery_index ? _T_257_199_0 : _GEN_1820;
  wire  _GEN_1825 = 8'hc7 == io_fetchQuery_index ? _T_257_199_1 : _GEN_1821;
  wire  _GEN_1826 = 8'hc7 == io_fetchQuery_index ? _T_257_199_2 : _GEN_1822;
  wire  _GEN_1827 = 8'hc7 == io_fetchQuery_index ? _T_257_199_3 : _GEN_1823;
  wire  _GEN_1828 = 8'hc8 == io_fetchQuery_index ? _T_257_200_0 : _GEN_1824;
  wire  _GEN_1829 = 8'hc8 == io_fetchQuery_index ? _T_257_200_1 : _GEN_1825;
  wire  _GEN_1830 = 8'hc8 == io_fetchQuery_index ? _T_257_200_2 : _GEN_1826;
  wire  _GEN_1831 = 8'hc8 == io_fetchQuery_index ? _T_257_200_3 : _GEN_1827;
  wire  _GEN_1832 = 8'hc9 == io_fetchQuery_index ? _T_257_201_0 : _GEN_1828;
  wire  _GEN_1833 = 8'hc9 == io_fetchQuery_index ? _T_257_201_1 : _GEN_1829;
  wire  _GEN_1834 = 8'hc9 == io_fetchQuery_index ? _T_257_201_2 : _GEN_1830;
  wire  _GEN_1835 = 8'hc9 == io_fetchQuery_index ? _T_257_201_3 : _GEN_1831;
  wire  _GEN_1836 = 8'hca == io_fetchQuery_index ? _T_257_202_0 : _GEN_1832;
  wire  _GEN_1837 = 8'hca == io_fetchQuery_index ? _T_257_202_1 : _GEN_1833;
  wire  _GEN_1838 = 8'hca == io_fetchQuery_index ? _T_257_202_2 : _GEN_1834;
  wire  _GEN_1839 = 8'hca == io_fetchQuery_index ? _T_257_202_3 : _GEN_1835;
  wire  _GEN_1840 = 8'hcb == io_fetchQuery_index ? _T_257_203_0 : _GEN_1836;
  wire  _GEN_1841 = 8'hcb == io_fetchQuery_index ? _T_257_203_1 : _GEN_1837;
  wire  _GEN_1842 = 8'hcb == io_fetchQuery_index ? _T_257_203_2 : _GEN_1838;
  wire  _GEN_1843 = 8'hcb == io_fetchQuery_index ? _T_257_203_3 : _GEN_1839;
  wire  _GEN_1844 = 8'hcc == io_fetchQuery_index ? _T_257_204_0 : _GEN_1840;
  wire  _GEN_1845 = 8'hcc == io_fetchQuery_index ? _T_257_204_1 : _GEN_1841;
  wire  _GEN_1846 = 8'hcc == io_fetchQuery_index ? _T_257_204_2 : _GEN_1842;
  wire  _GEN_1847 = 8'hcc == io_fetchQuery_index ? _T_257_204_3 : _GEN_1843;
  wire  _GEN_1848 = 8'hcd == io_fetchQuery_index ? _T_257_205_0 : _GEN_1844;
  wire  _GEN_1849 = 8'hcd == io_fetchQuery_index ? _T_257_205_1 : _GEN_1845;
  wire  _GEN_1850 = 8'hcd == io_fetchQuery_index ? _T_257_205_2 : _GEN_1846;
  wire  _GEN_1851 = 8'hcd == io_fetchQuery_index ? _T_257_205_3 : _GEN_1847;
  wire  _GEN_1852 = 8'hce == io_fetchQuery_index ? _T_257_206_0 : _GEN_1848;
  wire  _GEN_1853 = 8'hce == io_fetchQuery_index ? _T_257_206_1 : _GEN_1849;
  wire  _GEN_1854 = 8'hce == io_fetchQuery_index ? _T_257_206_2 : _GEN_1850;
  wire  _GEN_1855 = 8'hce == io_fetchQuery_index ? _T_257_206_3 : _GEN_1851;
  wire  _GEN_1856 = 8'hcf == io_fetchQuery_index ? _T_257_207_0 : _GEN_1852;
  wire  _GEN_1857 = 8'hcf == io_fetchQuery_index ? _T_257_207_1 : _GEN_1853;
  wire  _GEN_1858 = 8'hcf == io_fetchQuery_index ? _T_257_207_2 : _GEN_1854;
  wire  _GEN_1859 = 8'hcf == io_fetchQuery_index ? _T_257_207_3 : _GEN_1855;
  wire  _GEN_1860 = 8'hd0 == io_fetchQuery_index ? _T_257_208_0 : _GEN_1856;
  wire  _GEN_1861 = 8'hd0 == io_fetchQuery_index ? _T_257_208_1 : _GEN_1857;
  wire  _GEN_1862 = 8'hd0 == io_fetchQuery_index ? _T_257_208_2 : _GEN_1858;
  wire  _GEN_1863 = 8'hd0 == io_fetchQuery_index ? _T_257_208_3 : _GEN_1859;
  wire  _GEN_1864 = 8'hd1 == io_fetchQuery_index ? _T_257_209_0 : _GEN_1860;
  wire  _GEN_1865 = 8'hd1 == io_fetchQuery_index ? _T_257_209_1 : _GEN_1861;
  wire  _GEN_1866 = 8'hd1 == io_fetchQuery_index ? _T_257_209_2 : _GEN_1862;
  wire  _GEN_1867 = 8'hd1 == io_fetchQuery_index ? _T_257_209_3 : _GEN_1863;
  wire  _GEN_1868 = 8'hd2 == io_fetchQuery_index ? _T_257_210_0 : _GEN_1864;
  wire  _GEN_1869 = 8'hd2 == io_fetchQuery_index ? _T_257_210_1 : _GEN_1865;
  wire  _GEN_1870 = 8'hd2 == io_fetchQuery_index ? _T_257_210_2 : _GEN_1866;
  wire  _GEN_1871 = 8'hd2 == io_fetchQuery_index ? _T_257_210_3 : _GEN_1867;
  wire  _GEN_1872 = 8'hd3 == io_fetchQuery_index ? _T_257_211_0 : _GEN_1868;
  wire  _GEN_1873 = 8'hd3 == io_fetchQuery_index ? _T_257_211_1 : _GEN_1869;
  wire  _GEN_1874 = 8'hd3 == io_fetchQuery_index ? _T_257_211_2 : _GEN_1870;
  wire  _GEN_1875 = 8'hd3 == io_fetchQuery_index ? _T_257_211_3 : _GEN_1871;
  wire  _GEN_1876 = 8'hd4 == io_fetchQuery_index ? _T_257_212_0 : _GEN_1872;
  wire  _GEN_1877 = 8'hd4 == io_fetchQuery_index ? _T_257_212_1 : _GEN_1873;
  wire  _GEN_1878 = 8'hd4 == io_fetchQuery_index ? _T_257_212_2 : _GEN_1874;
  wire  _GEN_1879 = 8'hd4 == io_fetchQuery_index ? _T_257_212_3 : _GEN_1875;
  wire  _GEN_1880 = 8'hd5 == io_fetchQuery_index ? _T_257_213_0 : _GEN_1876;
  wire  _GEN_1881 = 8'hd5 == io_fetchQuery_index ? _T_257_213_1 : _GEN_1877;
  wire  _GEN_1882 = 8'hd5 == io_fetchQuery_index ? _T_257_213_2 : _GEN_1878;
  wire  _GEN_1883 = 8'hd5 == io_fetchQuery_index ? _T_257_213_3 : _GEN_1879;
  wire  _GEN_1884 = 8'hd6 == io_fetchQuery_index ? _T_257_214_0 : _GEN_1880;
  wire  _GEN_1885 = 8'hd6 == io_fetchQuery_index ? _T_257_214_1 : _GEN_1881;
  wire  _GEN_1886 = 8'hd6 == io_fetchQuery_index ? _T_257_214_2 : _GEN_1882;
  wire  _GEN_1887 = 8'hd6 == io_fetchQuery_index ? _T_257_214_3 : _GEN_1883;
  wire  _GEN_1888 = 8'hd7 == io_fetchQuery_index ? _T_257_215_0 : _GEN_1884;
  wire  _GEN_1889 = 8'hd7 == io_fetchQuery_index ? _T_257_215_1 : _GEN_1885;
  wire  _GEN_1890 = 8'hd7 == io_fetchQuery_index ? _T_257_215_2 : _GEN_1886;
  wire  _GEN_1891 = 8'hd7 == io_fetchQuery_index ? _T_257_215_3 : _GEN_1887;
  wire  _GEN_1892 = 8'hd8 == io_fetchQuery_index ? _T_257_216_0 : _GEN_1888;
  wire  _GEN_1893 = 8'hd8 == io_fetchQuery_index ? _T_257_216_1 : _GEN_1889;
  wire  _GEN_1894 = 8'hd8 == io_fetchQuery_index ? _T_257_216_2 : _GEN_1890;
  wire  _GEN_1895 = 8'hd8 == io_fetchQuery_index ? _T_257_216_3 : _GEN_1891;
  wire  _GEN_1896 = 8'hd9 == io_fetchQuery_index ? _T_257_217_0 : _GEN_1892;
  wire  _GEN_1897 = 8'hd9 == io_fetchQuery_index ? _T_257_217_1 : _GEN_1893;
  wire  _GEN_1898 = 8'hd9 == io_fetchQuery_index ? _T_257_217_2 : _GEN_1894;
  wire  _GEN_1899 = 8'hd9 == io_fetchQuery_index ? _T_257_217_3 : _GEN_1895;
  wire  _GEN_1900 = 8'hda == io_fetchQuery_index ? _T_257_218_0 : _GEN_1896;
  wire  _GEN_1901 = 8'hda == io_fetchQuery_index ? _T_257_218_1 : _GEN_1897;
  wire  _GEN_1902 = 8'hda == io_fetchQuery_index ? _T_257_218_2 : _GEN_1898;
  wire  _GEN_1903 = 8'hda == io_fetchQuery_index ? _T_257_218_3 : _GEN_1899;
  wire  _GEN_1904 = 8'hdb == io_fetchQuery_index ? _T_257_219_0 : _GEN_1900;
  wire  _GEN_1905 = 8'hdb == io_fetchQuery_index ? _T_257_219_1 : _GEN_1901;
  wire  _GEN_1906 = 8'hdb == io_fetchQuery_index ? _T_257_219_2 : _GEN_1902;
  wire  _GEN_1907 = 8'hdb == io_fetchQuery_index ? _T_257_219_3 : _GEN_1903;
  wire  _GEN_1908 = 8'hdc == io_fetchQuery_index ? _T_257_220_0 : _GEN_1904;
  wire  _GEN_1909 = 8'hdc == io_fetchQuery_index ? _T_257_220_1 : _GEN_1905;
  wire  _GEN_1910 = 8'hdc == io_fetchQuery_index ? _T_257_220_2 : _GEN_1906;
  wire  _GEN_1911 = 8'hdc == io_fetchQuery_index ? _T_257_220_3 : _GEN_1907;
  wire  _GEN_1912 = 8'hdd == io_fetchQuery_index ? _T_257_221_0 : _GEN_1908;
  wire  _GEN_1913 = 8'hdd == io_fetchQuery_index ? _T_257_221_1 : _GEN_1909;
  wire  _GEN_1914 = 8'hdd == io_fetchQuery_index ? _T_257_221_2 : _GEN_1910;
  wire  _GEN_1915 = 8'hdd == io_fetchQuery_index ? _T_257_221_3 : _GEN_1911;
  wire  _GEN_1916 = 8'hde == io_fetchQuery_index ? _T_257_222_0 : _GEN_1912;
  wire  _GEN_1917 = 8'hde == io_fetchQuery_index ? _T_257_222_1 : _GEN_1913;
  wire  _GEN_1918 = 8'hde == io_fetchQuery_index ? _T_257_222_2 : _GEN_1914;
  wire  _GEN_1919 = 8'hde == io_fetchQuery_index ? _T_257_222_3 : _GEN_1915;
  wire  _GEN_1920 = 8'hdf == io_fetchQuery_index ? _T_257_223_0 : _GEN_1916;
  wire  _GEN_1921 = 8'hdf == io_fetchQuery_index ? _T_257_223_1 : _GEN_1917;
  wire  _GEN_1922 = 8'hdf == io_fetchQuery_index ? _T_257_223_2 : _GEN_1918;
  wire  _GEN_1923 = 8'hdf == io_fetchQuery_index ? _T_257_223_3 : _GEN_1919;
  wire  _GEN_1924 = 8'he0 == io_fetchQuery_index ? _T_257_224_0 : _GEN_1920;
  wire  _GEN_1925 = 8'he0 == io_fetchQuery_index ? _T_257_224_1 : _GEN_1921;
  wire  _GEN_1926 = 8'he0 == io_fetchQuery_index ? _T_257_224_2 : _GEN_1922;
  wire  _GEN_1927 = 8'he0 == io_fetchQuery_index ? _T_257_224_3 : _GEN_1923;
  wire  _GEN_1928 = 8'he1 == io_fetchQuery_index ? _T_257_225_0 : _GEN_1924;
  wire  _GEN_1929 = 8'he1 == io_fetchQuery_index ? _T_257_225_1 : _GEN_1925;
  wire  _GEN_1930 = 8'he1 == io_fetchQuery_index ? _T_257_225_2 : _GEN_1926;
  wire  _GEN_1931 = 8'he1 == io_fetchQuery_index ? _T_257_225_3 : _GEN_1927;
  wire  _GEN_1932 = 8'he2 == io_fetchQuery_index ? _T_257_226_0 : _GEN_1928;
  wire  _GEN_1933 = 8'he2 == io_fetchQuery_index ? _T_257_226_1 : _GEN_1929;
  wire  _GEN_1934 = 8'he2 == io_fetchQuery_index ? _T_257_226_2 : _GEN_1930;
  wire  _GEN_1935 = 8'he2 == io_fetchQuery_index ? _T_257_226_3 : _GEN_1931;
  wire  _GEN_1936 = 8'he3 == io_fetchQuery_index ? _T_257_227_0 : _GEN_1932;
  wire  _GEN_1937 = 8'he3 == io_fetchQuery_index ? _T_257_227_1 : _GEN_1933;
  wire  _GEN_1938 = 8'he3 == io_fetchQuery_index ? _T_257_227_2 : _GEN_1934;
  wire  _GEN_1939 = 8'he3 == io_fetchQuery_index ? _T_257_227_3 : _GEN_1935;
  wire  _GEN_1940 = 8'he4 == io_fetchQuery_index ? _T_257_228_0 : _GEN_1936;
  wire  _GEN_1941 = 8'he4 == io_fetchQuery_index ? _T_257_228_1 : _GEN_1937;
  wire  _GEN_1942 = 8'he4 == io_fetchQuery_index ? _T_257_228_2 : _GEN_1938;
  wire  _GEN_1943 = 8'he4 == io_fetchQuery_index ? _T_257_228_3 : _GEN_1939;
  wire  _GEN_1944 = 8'he5 == io_fetchQuery_index ? _T_257_229_0 : _GEN_1940;
  wire  _GEN_1945 = 8'he5 == io_fetchQuery_index ? _T_257_229_1 : _GEN_1941;
  wire  _GEN_1946 = 8'he5 == io_fetchQuery_index ? _T_257_229_2 : _GEN_1942;
  wire  _GEN_1947 = 8'he5 == io_fetchQuery_index ? _T_257_229_3 : _GEN_1943;
  wire  _GEN_1948 = 8'he6 == io_fetchQuery_index ? _T_257_230_0 : _GEN_1944;
  wire  _GEN_1949 = 8'he6 == io_fetchQuery_index ? _T_257_230_1 : _GEN_1945;
  wire  _GEN_1950 = 8'he6 == io_fetchQuery_index ? _T_257_230_2 : _GEN_1946;
  wire  _GEN_1951 = 8'he6 == io_fetchQuery_index ? _T_257_230_3 : _GEN_1947;
  wire  _GEN_1952 = 8'he7 == io_fetchQuery_index ? _T_257_231_0 : _GEN_1948;
  wire  _GEN_1953 = 8'he7 == io_fetchQuery_index ? _T_257_231_1 : _GEN_1949;
  wire  _GEN_1954 = 8'he7 == io_fetchQuery_index ? _T_257_231_2 : _GEN_1950;
  wire  _GEN_1955 = 8'he7 == io_fetchQuery_index ? _T_257_231_3 : _GEN_1951;
  wire  _GEN_1956 = 8'he8 == io_fetchQuery_index ? _T_257_232_0 : _GEN_1952;
  wire  _GEN_1957 = 8'he8 == io_fetchQuery_index ? _T_257_232_1 : _GEN_1953;
  wire  _GEN_1958 = 8'he8 == io_fetchQuery_index ? _T_257_232_2 : _GEN_1954;
  wire  _GEN_1959 = 8'he8 == io_fetchQuery_index ? _T_257_232_3 : _GEN_1955;
  wire  _GEN_1960 = 8'he9 == io_fetchQuery_index ? _T_257_233_0 : _GEN_1956;
  wire  _GEN_1961 = 8'he9 == io_fetchQuery_index ? _T_257_233_1 : _GEN_1957;
  wire  _GEN_1962 = 8'he9 == io_fetchQuery_index ? _T_257_233_2 : _GEN_1958;
  wire  _GEN_1963 = 8'he9 == io_fetchQuery_index ? _T_257_233_3 : _GEN_1959;
  wire  _GEN_1964 = 8'hea == io_fetchQuery_index ? _T_257_234_0 : _GEN_1960;
  wire  _GEN_1965 = 8'hea == io_fetchQuery_index ? _T_257_234_1 : _GEN_1961;
  wire  _GEN_1966 = 8'hea == io_fetchQuery_index ? _T_257_234_2 : _GEN_1962;
  wire  _GEN_1967 = 8'hea == io_fetchQuery_index ? _T_257_234_3 : _GEN_1963;
  wire  _GEN_1968 = 8'heb == io_fetchQuery_index ? _T_257_235_0 : _GEN_1964;
  wire  _GEN_1969 = 8'heb == io_fetchQuery_index ? _T_257_235_1 : _GEN_1965;
  wire  _GEN_1970 = 8'heb == io_fetchQuery_index ? _T_257_235_2 : _GEN_1966;
  wire  _GEN_1971 = 8'heb == io_fetchQuery_index ? _T_257_235_3 : _GEN_1967;
  wire  _GEN_1972 = 8'hec == io_fetchQuery_index ? _T_257_236_0 : _GEN_1968;
  wire  _GEN_1973 = 8'hec == io_fetchQuery_index ? _T_257_236_1 : _GEN_1969;
  wire  _GEN_1974 = 8'hec == io_fetchQuery_index ? _T_257_236_2 : _GEN_1970;
  wire  _GEN_1975 = 8'hec == io_fetchQuery_index ? _T_257_236_3 : _GEN_1971;
  wire  _GEN_1976 = 8'hed == io_fetchQuery_index ? _T_257_237_0 : _GEN_1972;
  wire  _GEN_1977 = 8'hed == io_fetchQuery_index ? _T_257_237_1 : _GEN_1973;
  wire  _GEN_1978 = 8'hed == io_fetchQuery_index ? _T_257_237_2 : _GEN_1974;
  wire  _GEN_1979 = 8'hed == io_fetchQuery_index ? _T_257_237_3 : _GEN_1975;
  wire  _GEN_1980 = 8'hee == io_fetchQuery_index ? _T_257_238_0 : _GEN_1976;
  wire  _GEN_1981 = 8'hee == io_fetchQuery_index ? _T_257_238_1 : _GEN_1977;
  wire  _GEN_1982 = 8'hee == io_fetchQuery_index ? _T_257_238_2 : _GEN_1978;
  wire  _GEN_1983 = 8'hee == io_fetchQuery_index ? _T_257_238_3 : _GEN_1979;
  wire  _GEN_1984 = 8'hef == io_fetchQuery_index ? _T_257_239_0 : _GEN_1980;
  wire  _GEN_1985 = 8'hef == io_fetchQuery_index ? _T_257_239_1 : _GEN_1981;
  wire  _GEN_1986 = 8'hef == io_fetchQuery_index ? _T_257_239_2 : _GEN_1982;
  wire  _GEN_1987 = 8'hef == io_fetchQuery_index ? _T_257_239_3 : _GEN_1983;
  wire  _GEN_1988 = 8'hf0 == io_fetchQuery_index ? _T_257_240_0 : _GEN_1984;
  wire  _GEN_1989 = 8'hf0 == io_fetchQuery_index ? _T_257_240_1 : _GEN_1985;
  wire  _GEN_1990 = 8'hf0 == io_fetchQuery_index ? _T_257_240_2 : _GEN_1986;
  wire  _GEN_1991 = 8'hf0 == io_fetchQuery_index ? _T_257_240_3 : _GEN_1987;
  wire  _GEN_1992 = 8'hf1 == io_fetchQuery_index ? _T_257_241_0 : _GEN_1988;
  wire  _GEN_1993 = 8'hf1 == io_fetchQuery_index ? _T_257_241_1 : _GEN_1989;
  wire  _GEN_1994 = 8'hf1 == io_fetchQuery_index ? _T_257_241_2 : _GEN_1990;
  wire  _GEN_1995 = 8'hf1 == io_fetchQuery_index ? _T_257_241_3 : _GEN_1991;
  wire  _GEN_1996 = 8'hf2 == io_fetchQuery_index ? _T_257_242_0 : _GEN_1992;
  wire  _GEN_1997 = 8'hf2 == io_fetchQuery_index ? _T_257_242_1 : _GEN_1993;
  wire  _GEN_1998 = 8'hf2 == io_fetchQuery_index ? _T_257_242_2 : _GEN_1994;
  wire  _GEN_1999 = 8'hf2 == io_fetchQuery_index ? _T_257_242_3 : _GEN_1995;
  wire  _GEN_2000 = 8'hf3 == io_fetchQuery_index ? _T_257_243_0 : _GEN_1996;
  wire  _GEN_2001 = 8'hf3 == io_fetchQuery_index ? _T_257_243_1 : _GEN_1997;
  wire  _GEN_2002 = 8'hf3 == io_fetchQuery_index ? _T_257_243_2 : _GEN_1998;
  wire  _GEN_2003 = 8'hf3 == io_fetchQuery_index ? _T_257_243_3 : _GEN_1999;
  wire  _GEN_2004 = 8'hf4 == io_fetchQuery_index ? _T_257_244_0 : _GEN_2000;
  wire  _GEN_2005 = 8'hf4 == io_fetchQuery_index ? _T_257_244_1 : _GEN_2001;
  wire  _GEN_2006 = 8'hf4 == io_fetchQuery_index ? _T_257_244_2 : _GEN_2002;
  wire  _GEN_2007 = 8'hf4 == io_fetchQuery_index ? _T_257_244_3 : _GEN_2003;
  wire  _GEN_2008 = 8'hf5 == io_fetchQuery_index ? _T_257_245_0 : _GEN_2004;
  wire  _GEN_2009 = 8'hf5 == io_fetchQuery_index ? _T_257_245_1 : _GEN_2005;
  wire  _GEN_2010 = 8'hf5 == io_fetchQuery_index ? _T_257_245_2 : _GEN_2006;
  wire  _GEN_2011 = 8'hf5 == io_fetchQuery_index ? _T_257_245_3 : _GEN_2007;
  wire  _GEN_2012 = 8'hf6 == io_fetchQuery_index ? _T_257_246_0 : _GEN_2008;
  wire  _GEN_2013 = 8'hf6 == io_fetchQuery_index ? _T_257_246_1 : _GEN_2009;
  wire  _GEN_2014 = 8'hf6 == io_fetchQuery_index ? _T_257_246_2 : _GEN_2010;
  wire  _GEN_2015 = 8'hf6 == io_fetchQuery_index ? _T_257_246_3 : _GEN_2011;
  wire  _GEN_2016 = 8'hf7 == io_fetchQuery_index ? _T_257_247_0 : _GEN_2012;
  wire  _GEN_2017 = 8'hf7 == io_fetchQuery_index ? _T_257_247_1 : _GEN_2013;
  wire  _GEN_2018 = 8'hf7 == io_fetchQuery_index ? _T_257_247_2 : _GEN_2014;
  wire  _GEN_2019 = 8'hf7 == io_fetchQuery_index ? _T_257_247_3 : _GEN_2015;
  wire  _GEN_2020 = 8'hf8 == io_fetchQuery_index ? _T_257_248_0 : _GEN_2016;
  wire  _GEN_2021 = 8'hf8 == io_fetchQuery_index ? _T_257_248_1 : _GEN_2017;
  wire  _GEN_2022 = 8'hf8 == io_fetchQuery_index ? _T_257_248_2 : _GEN_2018;
  wire  _GEN_2023 = 8'hf8 == io_fetchQuery_index ? _T_257_248_3 : _GEN_2019;
  wire  _GEN_2024 = 8'hf9 == io_fetchQuery_index ? _T_257_249_0 : _GEN_2020;
  wire  _GEN_2025 = 8'hf9 == io_fetchQuery_index ? _T_257_249_1 : _GEN_2021;
  wire  _GEN_2026 = 8'hf9 == io_fetchQuery_index ? _T_257_249_2 : _GEN_2022;
  wire  _GEN_2027 = 8'hf9 == io_fetchQuery_index ? _T_257_249_3 : _GEN_2023;
  wire  _GEN_2028 = 8'hfa == io_fetchQuery_index ? _T_257_250_0 : _GEN_2024;
  wire  _GEN_2029 = 8'hfa == io_fetchQuery_index ? _T_257_250_1 : _GEN_2025;
  wire  _GEN_2030 = 8'hfa == io_fetchQuery_index ? _T_257_250_2 : _GEN_2026;
  wire  _GEN_2031 = 8'hfa == io_fetchQuery_index ? _T_257_250_3 : _GEN_2027;
  wire  _GEN_2032 = 8'hfb == io_fetchQuery_index ? _T_257_251_0 : _GEN_2028;
  wire  _GEN_2033 = 8'hfb == io_fetchQuery_index ? _T_257_251_1 : _GEN_2029;
  wire  _GEN_2034 = 8'hfb == io_fetchQuery_index ? _T_257_251_2 : _GEN_2030;
  wire  _GEN_2035 = 8'hfb == io_fetchQuery_index ? _T_257_251_3 : _GEN_2031;
  wire  _GEN_2036 = 8'hfc == io_fetchQuery_index ? _T_257_252_0 : _GEN_2032;
  wire  _GEN_2037 = 8'hfc == io_fetchQuery_index ? _T_257_252_1 : _GEN_2033;
  wire  _GEN_2038 = 8'hfc == io_fetchQuery_index ? _T_257_252_2 : _GEN_2034;
  wire  _GEN_2039 = 8'hfc == io_fetchQuery_index ? _T_257_252_3 : _GEN_2035;
  wire  _GEN_2040 = 8'hfd == io_fetchQuery_index ? _T_257_253_0 : _GEN_2036;
  wire  _GEN_2041 = 8'hfd == io_fetchQuery_index ? _T_257_253_1 : _GEN_2037;
  wire  _GEN_2042 = 8'hfd == io_fetchQuery_index ? _T_257_253_2 : _GEN_2038;
  wire  _GEN_2043 = 8'hfd == io_fetchQuery_index ? _T_257_253_3 : _GEN_2039;
  wire  _GEN_2044 = 8'hfe == io_fetchQuery_index ? _T_257_254_0 : _GEN_2040;
  wire  _GEN_2045 = 8'hfe == io_fetchQuery_index ? _T_257_254_1 : _GEN_2041;
  wire  _GEN_2046 = 8'hfe == io_fetchQuery_index ? _T_257_254_2 : _GEN_2042;
  wire  _GEN_2047 = 8'hfe == io_fetchQuery_index ? _T_257_254_3 : _GEN_2043;
  wire  _GEN_2048 = 8'hff == io_fetchQuery_index ? _T_257_255_0 : _GEN_2044;
  wire  _GEN_2049 = 8'hff == io_fetchQuery_index ? _T_257_255_1 : _GEN_2045;
  wire  _GEN_2050 = 8'hff == io_fetchQuery_index ? _T_257_255_2 : _GEN_2046;
  wire  _GEN_2051 = 8'hff == io_fetchQuery_index ? _T_257_255_3 : _GEN_2047;
  wire  _GEN_4108 = 2'h0 == comparator_io_bankHitWay_bits; // @[PLRUMRUNM.scala 25:21]
  wire  _GEN_2052 = _GEN_4108 | _GEN_2048; // @[PLRUMRUNM.scala 25:21]
  wire  _GEN_4109 = 2'h1 == comparator_io_bankHitWay_bits; // @[PLRUMRUNM.scala 25:21]
  wire  _GEN_2053 = _GEN_4109 | _GEN_2049; // @[PLRUMRUNM.scala 25:21]
  wire  _GEN_4110 = 2'h2 == comparator_io_bankHitWay_bits; // @[PLRUMRUNM.scala 25:21]
  wire  _GEN_2054 = _GEN_4110 | _GEN_2050; // @[PLRUMRUNM.scala 25:21]
  wire  _GEN_4111 = 2'h3 == comparator_io_bankHitWay_bits; // @[PLRUMRUNM.scala 25:21]
  wire  _GEN_2055 = _GEN_4111 | _GEN_2051; // @[PLRUMRUNM.scala 25:21]
  wire [3:0] _T_299 = {_GEN_2055,_GEN_2054,_GEN_2053,_GEN_2052}; // @[PLRUMRUNM.scala 28:37]
  wire  _T_300 = &_T_299; // @[PLRUMRUNM.scala 28:44]
  wire  _T_301_0 = _T_300 ? _GEN_4108 : _GEN_2052; // @[PLRUMRUNM.scala 28:25]
  wire  _T_301_1 = _T_300 ? _GEN_4109 : _GEN_2053; // @[PLRUMRUNM.scala 28:25]
  wire  _T_301_2 = _T_300 ? _GEN_4110 : _GEN_2054; // @[PLRUMRUNM.scala 28:25]
  wire  _T_301_3 = _T_300 ? _GEN_4111 : _GEN_2055; // @[PLRUMRUNM.scala 28:25]
  MSHR mshr ( // @[QueryTop.scala 37:28]
    .clock(mshr_clock),
    .reset(mshr_reset),
    .io_missAddr_ready(mshr_io_missAddr_ready),
    .io_missAddr_valid(mshr_io_missAddr_valid),
    .io_missAddr_bits_tag(mshr_io_missAddr_bits_tag),
    .io_missAddr_bits_index(mshr_io_missAddr_bits_index),
    .io_missAddr_bits_bankIndex(mshr_io_missAddr_bits_bankIndex),
    .io_readyForWB(mshr_io_readyForWB),
    .io_writeBack(mshr_io_writeBack),
    .io_mshrInfo_tag(mshr_io_mshrInfo_tag),
    .io_mshrInfo_index(mshr_io_mshrInfo_index),
    .io_mshrInfo_bankIndex(mshr_io_mshrInfo_bankIndex)
  );
  MissComparator comparator ( // @[QueryTop.scala 38:28]
    .io_tagValid_0_tag(comparator_io_tagValid_0_tag),
    .io_tagValid_0_valid(comparator_io_tagValid_0_valid),
    .io_tagValid_1_tag(comparator_io_tagValid_1_tag),
    .io_tagValid_1_valid(comparator_io_tagValid_1_valid),
    .io_tagValid_2_tag(comparator_io_tagValid_2_tag),
    .io_tagValid_2_valid(comparator_io_tagValid_2_valid),
    .io_tagValid_3_tag(comparator_io_tagValid_3_tag),
    .io_tagValid_3_valid(comparator_io_tagValid_3_valid),
    .io_phyTag(comparator_io_phyTag),
    .io_index(comparator_io_index),
    .io_mshr_bits_tag(comparator_io_mshr_bits_tag),
    .io_mshr_bits_index(comparator_io_mshr_bits_index),
    .io_refillBufferValid(comparator_io_refillBufferValid),
    .io_bankHitWay_valid(comparator_io_bankHitWay_valid),
    .io_bankHitWay_bits(comparator_io_bankHitWay_bits),
    .io_hitInRefillBuffer(comparator_io_hitInRefillBuffer)
  );
  AXIReadPort axi ( // @[QueryTop.scala 39:28]
    .clock(axi_clock),
    .reset(axi_reset),
    .io_axi_ar_ready(axi_io_axi_ar_ready),
    .io_axi_ar_valid(axi_io_axi_ar_valid),
    .io_axi_ar_bits_addr(axi_io_axi_ar_bits_addr),
    .io_axi_r_ready(axi_io_axi_r_ready),
    .io_axi_r_valid(axi_io_axi_r_valid),
    .io_axi_r_bits_data(axi_io_axi_r_bits_data),
    .io_axi_r_bits_last(axi_io_axi_r_bits_last),
    .io_addrReq_valid(axi_io_addrReq_valid),
    .io_addrReq_bits(axi_io_addrReq_bits),
    .io_transferData_valid(axi_io_transferData_valid),
    .io_transferData_bits(axi_io_transferData_bits),
    .io_finishTransfer(axi_io_finishTransfer)
  );
  ReFillBuffer refillBuffer ( // @[QueryTop.scala 40:28]
    .clock(refillBuffer_clock),
    .reset(refillBuffer_reset),
    .io_addr_valid(refillBuffer_io_addr_valid),
    .io_addr_bits(refillBuffer_io_addr_bits),
    .io_inputData_valid(refillBuffer_io_inputData_valid),
    .io_inputData_bits(refillBuffer_io_inputData_bits),
    .io_finish(refillBuffer_io_finish),
    .io_queryResult_valid(refillBuffer_io_queryResult_valid),
    .io_queryResult_bits(refillBuffer_io_queryResult_bits),
    .io_allData_0(refillBuffer_io_allData_0),
    .io_allData_1(refillBuffer_io_allData_1)
  );
  ReadHolder readHolder ( // @[QueryTop.scala 42:28]
    .clock(readHolder_clock),
    .reset(readHolder_reset),
    .io_input_valid(readHolder_io_input_valid),
    .io_input_bits(readHolder_io_input_bits),
    .io_output_valid(readHolder_io_output_valid),
    .io_output_bits(readHolder_io_output_bits)
  );
  assign io_ready = _T_264 | passThrough; // @[QueryTop.scala 64:17]
  assign io_data_valid = queryHit & _T_262; // @[QueryTop.scala 65:17]
  assign io_data_bits = readHolder_io_output_valid ? readHolder_io_output_bits : _T_266; // @[QueryTop.scala 66:16]
  assign io_writeBundle_writeEnable = mshr_io_writeBack; // @[QueryTop.scala 76:30]
  assign io_writeBundle_writeWay = _T_273 ? 2'h3 : _T_275; // @[QueryTop.scala 77:30]
  assign io_writeBundle_writeIndex = mshr_io_mshrInfo_index; // @[QueryTop.scala 78:30]
  assign io_writeBundle_writeTag = mshr_io_mshrInfo_tag; // @[QueryTop.scala 79:30]
  assign io_writeBundle_writeData_0 = refillBuffer_io_allData_0; // @[QueryTop.scala 80:30]
  assign io_writeBundle_writeData_1 = refillBuffer_io_allData_1; // @[QueryTop.scala 80:30]
  assign io_axi_ar_valid = axi_io_axi_ar_valid; // @[QueryTop.scala 83:10]
  assign io_axi_ar_bits_addr = axi_io_axi_ar_bits_addr; // @[QueryTop.scala 83:10]
  assign io_axi_r_ready = axi_io_axi_r_ready; // @[QueryTop.scala 83:10]
  assign mshr_clock = clock;
  assign mshr_reset = reset;
  assign mshr_io_missAddr_valid = _T_291 & _T_262; // @[QueryTop.scala 120:35]
  assign mshr_io_missAddr_bits_tag = io_fetchQuery_phyTag; // @[QueryTop.scala 121:35]
  assign mshr_io_missAddr_bits_index = io_fetchQuery_index; // @[QueryTop.scala 122:35]
  assign mshr_io_missAddr_bits_bankIndex = io_fetchQuery_bankIndex; // @[QueryTop.scala 123:35]
  assign mshr_io_readyForWB = axi_io_finishTransfer; // @[QueryTop.scala 124:35]
  assign comparator_io_tagValid_0_tag = io_fetchQuery_tagValid_0_tag; // @[QueryTop.scala 85:35]
  assign comparator_io_tagValid_0_valid = io_fetchQuery_tagValid_0_valid; // @[QueryTop.scala 85:35]
  assign comparator_io_tagValid_1_tag = io_fetchQuery_tagValid_1_tag; // @[QueryTop.scala 85:35]
  assign comparator_io_tagValid_1_valid = io_fetchQuery_tagValid_1_valid; // @[QueryTop.scala 85:35]
  assign comparator_io_tagValid_2_tag = io_fetchQuery_tagValid_2_tag; // @[QueryTop.scala 85:35]
  assign comparator_io_tagValid_2_valid = io_fetchQuery_tagValid_2_valid; // @[QueryTop.scala 85:35]
  assign comparator_io_tagValid_3_tag = io_fetchQuery_tagValid_3_tag; // @[QueryTop.scala 85:35]
  assign comparator_io_tagValid_3_valid = io_fetchQuery_tagValid_3_valid; // @[QueryTop.scala 85:35]
  assign comparator_io_phyTag = io_fetchQuery_phyTag; // @[QueryTop.scala 86:35]
  assign comparator_io_index = io_fetchQuery_index; // @[QueryTop.scala 87:35]
  assign comparator_io_mshr_bits_tag = mshr_io_mshrInfo_tag; // @[QueryTop.scala 88:35]
  assign comparator_io_mshr_bits_index = mshr_io_mshrInfo_index; // @[QueryTop.scala 88:35]
  assign comparator_io_refillBufferValid = refillBuffer_io_queryResult_valid; // @[QueryTop.scala 91:35]
  assign axi_clock = clock;
  assign axi_reset = reset;
  assign axi_io_axi_ar_ready = io_axi_ar_ready; // @[QueryTop.scala 83:10]
  assign axi_io_axi_r_valid = io_axi_r_valid; // @[QueryTop.scala 83:10]
  assign axi_io_axi_r_bits_data = io_axi_r_bits_data; // @[QueryTop.scala 83:10]
  assign axi_io_axi_r_bits_last = io_axi_r_bits_last; // @[QueryTop.scala 83:10]
  assign axi_io_addrReq_valid = mshr_io_missAddr_ready & mshr_io_missAddr_valid; // @[QueryTop.scala 117:24]
  assign axi_io_addrReq_bits = {{1'd0}, _T_290}; // @[QueryTop.scala 107:23]
  assign refillBuffer_clock = clock;
  assign refillBuffer_reset = reset;
  assign refillBuffer_io_addr_valid = mshr_io_missAddr_ready & mshr_io_missAddr_valid; // @[QueryTop.scala 93:30]
  assign refillBuffer_io_addr_bits = io_fetchQuery_bankIndex; // @[QueryTop.scala 94:30]
  assign refillBuffer_io_inputData_valid = axi_io_transferData_valid; // @[QueryTop.scala 95:30]
  assign refillBuffer_io_inputData_bits = axi_io_transferData_bits; // @[QueryTop.scala 95:30]
  assign refillBuffer_io_finish = axi_io_finishTransfer; // @[QueryTop.scala 96:30]
  assign readHolder_clock = clock;
  assign readHolder_reset = reset;
  assign readHolder_io_input_valid = validData & _T_278; // @[QueryTop.scala 98:29]
  assign readHolder_io_input_bits = comparator_io_hitInRefillBuffer ? refillBuffer_io_queryResult_bits : _T_282; // @[QueryTop.scala 99:28]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_257_0_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  _T_257_0_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  _T_257_0_2 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  _T_257_0_3 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  _T_257_1_0 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  _T_257_1_1 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  _T_257_1_2 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  _T_257_1_3 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  _T_257_2_0 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  _T_257_2_1 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  _T_257_2_2 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  _T_257_2_3 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  _T_257_3_0 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  _T_257_3_1 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  _T_257_3_2 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  _T_257_3_3 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  _T_257_4_0 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  _T_257_4_1 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  _T_257_4_2 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  _T_257_4_3 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  _T_257_5_0 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  _T_257_5_1 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  _T_257_5_2 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  _T_257_5_3 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  _T_257_6_0 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  _T_257_6_1 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  _T_257_6_2 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  _T_257_6_3 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  _T_257_7_0 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  _T_257_7_1 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  _T_257_7_2 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  _T_257_7_3 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  _T_257_8_0 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  _T_257_8_1 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  _T_257_8_2 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  _T_257_8_3 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  _T_257_9_0 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  _T_257_9_1 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  _T_257_9_2 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  _T_257_9_3 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  _T_257_10_0 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  _T_257_10_1 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  _T_257_10_2 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  _T_257_10_3 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  _T_257_11_0 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  _T_257_11_1 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  _T_257_11_2 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  _T_257_11_3 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  _T_257_12_0 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  _T_257_12_1 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  _T_257_12_2 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  _T_257_12_3 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  _T_257_13_0 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  _T_257_13_1 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  _T_257_13_2 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  _T_257_13_3 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  _T_257_14_0 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  _T_257_14_1 = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  _T_257_14_2 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  _T_257_14_3 = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  _T_257_15_0 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  _T_257_15_1 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  _T_257_15_2 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  _T_257_15_3 = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  _T_257_16_0 = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  _T_257_16_1 = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  _T_257_16_2 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  _T_257_16_3 = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  _T_257_17_0 = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  _T_257_17_1 = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  _T_257_17_2 = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  _T_257_17_3 = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  _T_257_18_0 = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  _T_257_18_1 = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  _T_257_18_2 = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  _T_257_18_3 = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  _T_257_19_0 = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  _T_257_19_1 = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  _T_257_19_2 = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  _T_257_19_3 = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  _T_257_20_0 = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  _T_257_20_1 = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  _T_257_20_2 = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  _T_257_20_3 = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  _T_257_21_0 = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  _T_257_21_1 = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  _T_257_21_2 = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  _T_257_21_3 = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  _T_257_22_0 = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  _T_257_22_1 = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  _T_257_22_2 = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  _T_257_22_3 = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  _T_257_23_0 = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  _T_257_23_1 = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  _T_257_23_2 = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  _T_257_23_3 = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  _T_257_24_0 = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  _T_257_24_1 = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  _T_257_24_2 = _RAND_98[0:0];
  _RAND_99 = {1{`RANDOM}};
  _T_257_24_3 = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  _T_257_25_0 = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  _T_257_25_1 = _RAND_101[0:0];
  _RAND_102 = {1{`RANDOM}};
  _T_257_25_2 = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  _T_257_25_3 = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  _T_257_26_0 = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  _T_257_26_1 = _RAND_105[0:0];
  _RAND_106 = {1{`RANDOM}};
  _T_257_26_2 = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  _T_257_26_3 = _RAND_107[0:0];
  _RAND_108 = {1{`RANDOM}};
  _T_257_27_0 = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  _T_257_27_1 = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  _T_257_27_2 = _RAND_110[0:0];
  _RAND_111 = {1{`RANDOM}};
  _T_257_27_3 = _RAND_111[0:0];
  _RAND_112 = {1{`RANDOM}};
  _T_257_28_0 = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  _T_257_28_1 = _RAND_113[0:0];
  _RAND_114 = {1{`RANDOM}};
  _T_257_28_2 = _RAND_114[0:0];
  _RAND_115 = {1{`RANDOM}};
  _T_257_28_3 = _RAND_115[0:0];
  _RAND_116 = {1{`RANDOM}};
  _T_257_29_0 = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  _T_257_29_1 = _RAND_117[0:0];
  _RAND_118 = {1{`RANDOM}};
  _T_257_29_2 = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  _T_257_29_3 = _RAND_119[0:0];
  _RAND_120 = {1{`RANDOM}};
  _T_257_30_0 = _RAND_120[0:0];
  _RAND_121 = {1{`RANDOM}};
  _T_257_30_1 = _RAND_121[0:0];
  _RAND_122 = {1{`RANDOM}};
  _T_257_30_2 = _RAND_122[0:0];
  _RAND_123 = {1{`RANDOM}};
  _T_257_30_3 = _RAND_123[0:0];
  _RAND_124 = {1{`RANDOM}};
  _T_257_31_0 = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  _T_257_31_1 = _RAND_125[0:0];
  _RAND_126 = {1{`RANDOM}};
  _T_257_31_2 = _RAND_126[0:0];
  _RAND_127 = {1{`RANDOM}};
  _T_257_31_3 = _RAND_127[0:0];
  _RAND_128 = {1{`RANDOM}};
  _T_257_32_0 = _RAND_128[0:0];
  _RAND_129 = {1{`RANDOM}};
  _T_257_32_1 = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  _T_257_32_2 = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  _T_257_32_3 = _RAND_131[0:0];
  _RAND_132 = {1{`RANDOM}};
  _T_257_33_0 = _RAND_132[0:0];
  _RAND_133 = {1{`RANDOM}};
  _T_257_33_1 = _RAND_133[0:0];
  _RAND_134 = {1{`RANDOM}};
  _T_257_33_2 = _RAND_134[0:0];
  _RAND_135 = {1{`RANDOM}};
  _T_257_33_3 = _RAND_135[0:0];
  _RAND_136 = {1{`RANDOM}};
  _T_257_34_0 = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  _T_257_34_1 = _RAND_137[0:0];
  _RAND_138 = {1{`RANDOM}};
  _T_257_34_2 = _RAND_138[0:0];
  _RAND_139 = {1{`RANDOM}};
  _T_257_34_3 = _RAND_139[0:0];
  _RAND_140 = {1{`RANDOM}};
  _T_257_35_0 = _RAND_140[0:0];
  _RAND_141 = {1{`RANDOM}};
  _T_257_35_1 = _RAND_141[0:0];
  _RAND_142 = {1{`RANDOM}};
  _T_257_35_2 = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  _T_257_35_3 = _RAND_143[0:0];
  _RAND_144 = {1{`RANDOM}};
  _T_257_36_0 = _RAND_144[0:0];
  _RAND_145 = {1{`RANDOM}};
  _T_257_36_1 = _RAND_145[0:0];
  _RAND_146 = {1{`RANDOM}};
  _T_257_36_2 = _RAND_146[0:0];
  _RAND_147 = {1{`RANDOM}};
  _T_257_36_3 = _RAND_147[0:0];
  _RAND_148 = {1{`RANDOM}};
  _T_257_37_0 = _RAND_148[0:0];
  _RAND_149 = {1{`RANDOM}};
  _T_257_37_1 = _RAND_149[0:0];
  _RAND_150 = {1{`RANDOM}};
  _T_257_37_2 = _RAND_150[0:0];
  _RAND_151 = {1{`RANDOM}};
  _T_257_37_3 = _RAND_151[0:0];
  _RAND_152 = {1{`RANDOM}};
  _T_257_38_0 = _RAND_152[0:0];
  _RAND_153 = {1{`RANDOM}};
  _T_257_38_1 = _RAND_153[0:0];
  _RAND_154 = {1{`RANDOM}};
  _T_257_38_2 = _RAND_154[0:0];
  _RAND_155 = {1{`RANDOM}};
  _T_257_38_3 = _RAND_155[0:0];
  _RAND_156 = {1{`RANDOM}};
  _T_257_39_0 = _RAND_156[0:0];
  _RAND_157 = {1{`RANDOM}};
  _T_257_39_1 = _RAND_157[0:0];
  _RAND_158 = {1{`RANDOM}};
  _T_257_39_2 = _RAND_158[0:0];
  _RAND_159 = {1{`RANDOM}};
  _T_257_39_3 = _RAND_159[0:0];
  _RAND_160 = {1{`RANDOM}};
  _T_257_40_0 = _RAND_160[0:0];
  _RAND_161 = {1{`RANDOM}};
  _T_257_40_1 = _RAND_161[0:0];
  _RAND_162 = {1{`RANDOM}};
  _T_257_40_2 = _RAND_162[0:0];
  _RAND_163 = {1{`RANDOM}};
  _T_257_40_3 = _RAND_163[0:0];
  _RAND_164 = {1{`RANDOM}};
  _T_257_41_0 = _RAND_164[0:0];
  _RAND_165 = {1{`RANDOM}};
  _T_257_41_1 = _RAND_165[0:0];
  _RAND_166 = {1{`RANDOM}};
  _T_257_41_2 = _RAND_166[0:0];
  _RAND_167 = {1{`RANDOM}};
  _T_257_41_3 = _RAND_167[0:0];
  _RAND_168 = {1{`RANDOM}};
  _T_257_42_0 = _RAND_168[0:0];
  _RAND_169 = {1{`RANDOM}};
  _T_257_42_1 = _RAND_169[0:0];
  _RAND_170 = {1{`RANDOM}};
  _T_257_42_2 = _RAND_170[0:0];
  _RAND_171 = {1{`RANDOM}};
  _T_257_42_3 = _RAND_171[0:0];
  _RAND_172 = {1{`RANDOM}};
  _T_257_43_0 = _RAND_172[0:0];
  _RAND_173 = {1{`RANDOM}};
  _T_257_43_1 = _RAND_173[0:0];
  _RAND_174 = {1{`RANDOM}};
  _T_257_43_2 = _RAND_174[0:0];
  _RAND_175 = {1{`RANDOM}};
  _T_257_43_3 = _RAND_175[0:0];
  _RAND_176 = {1{`RANDOM}};
  _T_257_44_0 = _RAND_176[0:0];
  _RAND_177 = {1{`RANDOM}};
  _T_257_44_1 = _RAND_177[0:0];
  _RAND_178 = {1{`RANDOM}};
  _T_257_44_2 = _RAND_178[0:0];
  _RAND_179 = {1{`RANDOM}};
  _T_257_44_3 = _RAND_179[0:0];
  _RAND_180 = {1{`RANDOM}};
  _T_257_45_0 = _RAND_180[0:0];
  _RAND_181 = {1{`RANDOM}};
  _T_257_45_1 = _RAND_181[0:0];
  _RAND_182 = {1{`RANDOM}};
  _T_257_45_2 = _RAND_182[0:0];
  _RAND_183 = {1{`RANDOM}};
  _T_257_45_3 = _RAND_183[0:0];
  _RAND_184 = {1{`RANDOM}};
  _T_257_46_0 = _RAND_184[0:0];
  _RAND_185 = {1{`RANDOM}};
  _T_257_46_1 = _RAND_185[0:0];
  _RAND_186 = {1{`RANDOM}};
  _T_257_46_2 = _RAND_186[0:0];
  _RAND_187 = {1{`RANDOM}};
  _T_257_46_3 = _RAND_187[0:0];
  _RAND_188 = {1{`RANDOM}};
  _T_257_47_0 = _RAND_188[0:0];
  _RAND_189 = {1{`RANDOM}};
  _T_257_47_1 = _RAND_189[0:0];
  _RAND_190 = {1{`RANDOM}};
  _T_257_47_2 = _RAND_190[0:0];
  _RAND_191 = {1{`RANDOM}};
  _T_257_47_3 = _RAND_191[0:0];
  _RAND_192 = {1{`RANDOM}};
  _T_257_48_0 = _RAND_192[0:0];
  _RAND_193 = {1{`RANDOM}};
  _T_257_48_1 = _RAND_193[0:0];
  _RAND_194 = {1{`RANDOM}};
  _T_257_48_2 = _RAND_194[0:0];
  _RAND_195 = {1{`RANDOM}};
  _T_257_48_3 = _RAND_195[0:0];
  _RAND_196 = {1{`RANDOM}};
  _T_257_49_0 = _RAND_196[0:0];
  _RAND_197 = {1{`RANDOM}};
  _T_257_49_1 = _RAND_197[0:0];
  _RAND_198 = {1{`RANDOM}};
  _T_257_49_2 = _RAND_198[0:0];
  _RAND_199 = {1{`RANDOM}};
  _T_257_49_3 = _RAND_199[0:0];
  _RAND_200 = {1{`RANDOM}};
  _T_257_50_0 = _RAND_200[0:0];
  _RAND_201 = {1{`RANDOM}};
  _T_257_50_1 = _RAND_201[0:0];
  _RAND_202 = {1{`RANDOM}};
  _T_257_50_2 = _RAND_202[0:0];
  _RAND_203 = {1{`RANDOM}};
  _T_257_50_3 = _RAND_203[0:0];
  _RAND_204 = {1{`RANDOM}};
  _T_257_51_0 = _RAND_204[0:0];
  _RAND_205 = {1{`RANDOM}};
  _T_257_51_1 = _RAND_205[0:0];
  _RAND_206 = {1{`RANDOM}};
  _T_257_51_2 = _RAND_206[0:0];
  _RAND_207 = {1{`RANDOM}};
  _T_257_51_3 = _RAND_207[0:0];
  _RAND_208 = {1{`RANDOM}};
  _T_257_52_0 = _RAND_208[0:0];
  _RAND_209 = {1{`RANDOM}};
  _T_257_52_1 = _RAND_209[0:0];
  _RAND_210 = {1{`RANDOM}};
  _T_257_52_2 = _RAND_210[0:0];
  _RAND_211 = {1{`RANDOM}};
  _T_257_52_3 = _RAND_211[0:0];
  _RAND_212 = {1{`RANDOM}};
  _T_257_53_0 = _RAND_212[0:0];
  _RAND_213 = {1{`RANDOM}};
  _T_257_53_1 = _RAND_213[0:0];
  _RAND_214 = {1{`RANDOM}};
  _T_257_53_2 = _RAND_214[0:0];
  _RAND_215 = {1{`RANDOM}};
  _T_257_53_3 = _RAND_215[0:0];
  _RAND_216 = {1{`RANDOM}};
  _T_257_54_0 = _RAND_216[0:0];
  _RAND_217 = {1{`RANDOM}};
  _T_257_54_1 = _RAND_217[0:0];
  _RAND_218 = {1{`RANDOM}};
  _T_257_54_2 = _RAND_218[0:0];
  _RAND_219 = {1{`RANDOM}};
  _T_257_54_3 = _RAND_219[0:0];
  _RAND_220 = {1{`RANDOM}};
  _T_257_55_0 = _RAND_220[0:0];
  _RAND_221 = {1{`RANDOM}};
  _T_257_55_1 = _RAND_221[0:0];
  _RAND_222 = {1{`RANDOM}};
  _T_257_55_2 = _RAND_222[0:0];
  _RAND_223 = {1{`RANDOM}};
  _T_257_55_3 = _RAND_223[0:0];
  _RAND_224 = {1{`RANDOM}};
  _T_257_56_0 = _RAND_224[0:0];
  _RAND_225 = {1{`RANDOM}};
  _T_257_56_1 = _RAND_225[0:0];
  _RAND_226 = {1{`RANDOM}};
  _T_257_56_2 = _RAND_226[0:0];
  _RAND_227 = {1{`RANDOM}};
  _T_257_56_3 = _RAND_227[0:0];
  _RAND_228 = {1{`RANDOM}};
  _T_257_57_0 = _RAND_228[0:0];
  _RAND_229 = {1{`RANDOM}};
  _T_257_57_1 = _RAND_229[0:0];
  _RAND_230 = {1{`RANDOM}};
  _T_257_57_2 = _RAND_230[0:0];
  _RAND_231 = {1{`RANDOM}};
  _T_257_57_3 = _RAND_231[0:0];
  _RAND_232 = {1{`RANDOM}};
  _T_257_58_0 = _RAND_232[0:0];
  _RAND_233 = {1{`RANDOM}};
  _T_257_58_1 = _RAND_233[0:0];
  _RAND_234 = {1{`RANDOM}};
  _T_257_58_2 = _RAND_234[0:0];
  _RAND_235 = {1{`RANDOM}};
  _T_257_58_3 = _RAND_235[0:0];
  _RAND_236 = {1{`RANDOM}};
  _T_257_59_0 = _RAND_236[0:0];
  _RAND_237 = {1{`RANDOM}};
  _T_257_59_1 = _RAND_237[0:0];
  _RAND_238 = {1{`RANDOM}};
  _T_257_59_2 = _RAND_238[0:0];
  _RAND_239 = {1{`RANDOM}};
  _T_257_59_3 = _RAND_239[0:0];
  _RAND_240 = {1{`RANDOM}};
  _T_257_60_0 = _RAND_240[0:0];
  _RAND_241 = {1{`RANDOM}};
  _T_257_60_1 = _RAND_241[0:0];
  _RAND_242 = {1{`RANDOM}};
  _T_257_60_2 = _RAND_242[0:0];
  _RAND_243 = {1{`RANDOM}};
  _T_257_60_3 = _RAND_243[0:0];
  _RAND_244 = {1{`RANDOM}};
  _T_257_61_0 = _RAND_244[0:0];
  _RAND_245 = {1{`RANDOM}};
  _T_257_61_1 = _RAND_245[0:0];
  _RAND_246 = {1{`RANDOM}};
  _T_257_61_2 = _RAND_246[0:0];
  _RAND_247 = {1{`RANDOM}};
  _T_257_61_3 = _RAND_247[0:0];
  _RAND_248 = {1{`RANDOM}};
  _T_257_62_0 = _RAND_248[0:0];
  _RAND_249 = {1{`RANDOM}};
  _T_257_62_1 = _RAND_249[0:0];
  _RAND_250 = {1{`RANDOM}};
  _T_257_62_2 = _RAND_250[0:0];
  _RAND_251 = {1{`RANDOM}};
  _T_257_62_3 = _RAND_251[0:0];
  _RAND_252 = {1{`RANDOM}};
  _T_257_63_0 = _RAND_252[0:0];
  _RAND_253 = {1{`RANDOM}};
  _T_257_63_1 = _RAND_253[0:0];
  _RAND_254 = {1{`RANDOM}};
  _T_257_63_2 = _RAND_254[0:0];
  _RAND_255 = {1{`RANDOM}};
  _T_257_63_3 = _RAND_255[0:0];
  _RAND_256 = {1{`RANDOM}};
  _T_257_64_0 = _RAND_256[0:0];
  _RAND_257 = {1{`RANDOM}};
  _T_257_64_1 = _RAND_257[0:0];
  _RAND_258 = {1{`RANDOM}};
  _T_257_64_2 = _RAND_258[0:0];
  _RAND_259 = {1{`RANDOM}};
  _T_257_64_3 = _RAND_259[0:0];
  _RAND_260 = {1{`RANDOM}};
  _T_257_65_0 = _RAND_260[0:0];
  _RAND_261 = {1{`RANDOM}};
  _T_257_65_1 = _RAND_261[0:0];
  _RAND_262 = {1{`RANDOM}};
  _T_257_65_2 = _RAND_262[0:0];
  _RAND_263 = {1{`RANDOM}};
  _T_257_65_3 = _RAND_263[0:0];
  _RAND_264 = {1{`RANDOM}};
  _T_257_66_0 = _RAND_264[0:0];
  _RAND_265 = {1{`RANDOM}};
  _T_257_66_1 = _RAND_265[0:0];
  _RAND_266 = {1{`RANDOM}};
  _T_257_66_2 = _RAND_266[0:0];
  _RAND_267 = {1{`RANDOM}};
  _T_257_66_3 = _RAND_267[0:0];
  _RAND_268 = {1{`RANDOM}};
  _T_257_67_0 = _RAND_268[0:0];
  _RAND_269 = {1{`RANDOM}};
  _T_257_67_1 = _RAND_269[0:0];
  _RAND_270 = {1{`RANDOM}};
  _T_257_67_2 = _RAND_270[0:0];
  _RAND_271 = {1{`RANDOM}};
  _T_257_67_3 = _RAND_271[0:0];
  _RAND_272 = {1{`RANDOM}};
  _T_257_68_0 = _RAND_272[0:0];
  _RAND_273 = {1{`RANDOM}};
  _T_257_68_1 = _RAND_273[0:0];
  _RAND_274 = {1{`RANDOM}};
  _T_257_68_2 = _RAND_274[0:0];
  _RAND_275 = {1{`RANDOM}};
  _T_257_68_3 = _RAND_275[0:0];
  _RAND_276 = {1{`RANDOM}};
  _T_257_69_0 = _RAND_276[0:0];
  _RAND_277 = {1{`RANDOM}};
  _T_257_69_1 = _RAND_277[0:0];
  _RAND_278 = {1{`RANDOM}};
  _T_257_69_2 = _RAND_278[0:0];
  _RAND_279 = {1{`RANDOM}};
  _T_257_69_3 = _RAND_279[0:0];
  _RAND_280 = {1{`RANDOM}};
  _T_257_70_0 = _RAND_280[0:0];
  _RAND_281 = {1{`RANDOM}};
  _T_257_70_1 = _RAND_281[0:0];
  _RAND_282 = {1{`RANDOM}};
  _T_257_70_2 = _RAND_282[0:0];
  _RAND_283 = {1{`RANDOM}};
  _T_257_70_3 = _RAND_283[0:0];
  _RAND_284 = {1{`RANDOM}};
  _T_257_71_0 = _RAND_284[0:0];
  _RAND_285 = {1{`RANDOM}};
  _T_257_71_1 = _RAND_285[0:0];
  _RAND_286 = {1{`RANDOM}};
  _T_257_71_2 = _RAND_286[0:0];
  _RAND_287 = {1{`RANDOM}};
  _T_257_71_3 = _RAND_287[0:0];
  _RAND_288 = {1{`RANDOM}};
  _T_257_72_0 = _RAND_288[0:0];
  _RAND_289 = {1{`RANDOM}};
  _T_257_72_1 = _RAND_289[0:0];
  _RAND_290 = {1{`RANDOM}};
  _T_257_72_2 = _RAND_290[0:0];
  _RAND_291 = {1{`RANDOM}};
  _T_257_72_3 = _RAND_291[0:0];
  _RAND_292 = {1{`RANDOM}};
  _T_257_73_0 = _RAND_292[0:0];
  _RAND_293 = {1{`RANDOM}};
  _T_257_73_1 = _RAND_293[0:0];
  _RAND_294 = {1{`RANDOM}};
  _T_257_73_2 = _RAND_294[0:0];
  _RAND_295 = {1{`RANDOM}};
  _T_257_73_3 = _RAND_295[0:0];
  _RAND_296 = {1{`RANDOM}};
  _T_257_74_0 = _RAND_296[0:0];
  _RAND_297 = {1{`RANDOM}};
  _T_257_74_1 = _RAND_297[0:0];
  _RAND_298 = {1{`RANDOM}};
  _T_257_74_2 = _RAND_298[0:0];
  _RAND_299 = {1{`RANDOM}};
  _T_257_74_3 = _RAND_299[0:0];
  _RAND_300 = {1{`RANDOM}};
  _T_257_75_0 = _RAND_300[0:0];
  _RAND_301 = {1{`RANDOM}};
  _T_257_75_1 = _RAND_301[0:0];
  _RAND_302 = {1{`RANDOM}};
  _T_257_75_2 = _RAND_302[0:0];
  _RAND_303 = {1{`RANDOM}};
  _T_257_75_3 = _RAND_303[0:0];
  _RAND_304 = {1{`RANDOM}};
  _T_257_76_0 = _RAND_304[0:0];
  _RAND_305 = {1{`RANDOM}};
  _T_257_76_1 = _RAND_305[0:0];
  _RAND_306 = {1{`RANDOM}};
  _T_257_76_2 = _RAND_306[0:0];
  _RAND_307 = {1{`RANDOM}};
  _T_257_76_3 = _RAND_307[0:0];
  _RAND_308 = {1{`RANDOM}};
  _T_257_77_0 = _RAND_308[0:0];
  _RAND_309 = {1{`RANDOM}};
  _T_257_77_1 = _RAND_309[0:0];
  _RAND_310 = {1{`RANDOM}};
  _T_257_77_2 = _RAND_310[0:0];
  _RAND_311 = {1{`RANDOM}};
  _T_257_77_3 = _RAND_311[0:0];
  _RAND_312 = {1{`RANDOM}};
  _T_257_78_0 = _RAND_312[0:0];
  _RAND_313 = {1{`RANDOM}};
  _T_257_78_1 = _RAND_313[0:0];
  _RAND_314 = {1{`RANDOM}};
  _T_257_78_2 = _RAND_314[0:0];
  _RAND_315 = {1{`RANDOM}};
  _T_257_78_3 = _RAND_315[0:0];
  _RAND_316 = {1{`RANDOM}};
  _T_257_79_0 = _RAND_316[0:0];
  _RAND_317 = {1{`RANDOM}};
  _T_257_79_1 = _RAND_317[0:0];
  _RAND_318 = {1{`RANDOM}};
  _T_257_79_2 = _RAND_318[0:0];
  _RAND_319 = {1{`RANDOM}};
  _T_257_79_3 = _RAND_319[0:0];
  _RAND_320 = {1{`RANDOM}};
  _T_257_80_0 = _RAND_320[0:0];
  _RAND_321 = {1{`RANDOM}};
  _T_257_80_1 = _RAND_321[0:0];
  _RAND_322 = {1{`RANDOM}};
  _T_257_80_2 = _RAND_322[0:0];
  _RAND_323 = {1{`RANDOM}};
  _T_257_80_3 = _RAND_323[0:0];
  _RAND_324 = {1{`RANDOM}};
  _T_257_81_0 = _RAND_324[0:0];
  _RAND_325 = {1{`RANDOM}};
  _T_257_81_1 = _RAND_325[0:0];
  _RAND_326 = {1{`RANDOM}};
  _T_257_81_2 = _RAND_326[0:0];
  _RAND_327 = {1{`RANDOM}};
  _T_257_81_3 = _RAND_327[0:0];
  _RAND_328 = {1{`RANDOM}};
  _T_257_82_0 = _RAND_328[0:0];
  _RAND_329 = {1{`RANDOM}};
  _T_257_82_1 = _RAND_329[0:0];
  _RAND_330 = {1{`RANDOM}};
  _T_257_82_2 = _RAND_330[0:0];
  _RAND_331 = {1{`RANDOM}};
  _T_257_82_3 = _RAND_331[0:0];
  _RAND_332 = {1{`RANDOM}};
  _T_257_83_0 = _RAND_332[0:0];
  _RAND_333 = {1{`RANDOM}};
  _T_257_83_1 = _RAND_333[0:0];
  _RAND_334 = {1{`RANDOM}};
  _T_257_83_2 = _RAND_334[0:0];
  _RAND_335 = {1{`RANDOM}};
  _T_257_83_3 = _RAND_335[0:0];
  _RAND_336 = {1{`RANDOM}};
  _T_257_84_0 = _RAND_336[0:0];
  _RAND_337 = {1{`RANDOM}};
  _T_257_84_1 = _RAND_337[0:0];
  _RAND_338 = {1{`RANDOM}};
  _T_257_84_2 = _RAND_338[0:0];
  _RAND_339 = {1{`RANDOM}};
  _T_257_84_3 = _RAND_339[0:0];
  _RAND_340 = {1{`RANDOM}};
  _T_257_85_0 = _RAND_340[0:0];
  _RAND_341 = {1{`RANDOM}};
  _T_257_85_1 = _RAND_341[0:0];
  _RAND_342 = {1{`RANDOM}};
  _T_257_85_2 = _RAND_342[0:0];
  _RAND_343 = {1{`RANDOM}};
  _T_257_85_3 = _RAND_343[0:0];
  _RAND_344 = {1{`RANDOM}};
  _T_257_86_0 = _RAND_344[0:0];
  _RAND_345 = {1{`RANDOM}};
  _T_257_86_1 = _RAND_345[0:0];
  _RAND_346 = {1{`RANDOM}};
  _T_257_86_2 = _RAND_346[0:0];
  _RAND_347 = {1{`RANDOM}};
  _T_257_86_3 = _RAND_347[0:0];
  _RAND_348 = {1{`RANDOM}};
  _T_257_87_0 = _RAND_348[0:0];
  _RAND_349 = {1{`RANDOM}};
  _T_257_87_1 = _RAND_349[0:0];
  _RAND_350 = {1{`RANDOM}};
  _T_257_87_2 = _RAND_350[0:0];
  _RAND_351 = {1{`RANDOM}};
  _T_257_87_3 = _RAND_351[0:0];
  _RAND_352 = {1{`RANDOM}};
  _T_257_88_0 = _RAND_352[0:0];
  _RAND_353 = {1{`RANDOM}};
  _T_257_88_1 = _RAND_353[0:0];
  _RAND_354 = {1{`RANDOM}};
  _T_257_88_2 = _RAND_354[0:0];
  _RAND_355 = {1{`RANDOM}};
  _T_257_88_3 = _RAND_355[0:0];
  _RAND_356 = {1{`RANDOM}};
  _T_257_89_0 = _RAND_356[0:0];
  _RAND_357 = {1{`RANDOM}};
  _T_257_89_1 = _RAND_357[0:0];
  _RAND_358 = {1{`RANDOM}};
  _T_257_89_2 = _RAND_358[0:0];
  _RAND_359 = {1{`RANDOM}};
  _T_257_89_3 = _RAND_359[0:0];
  _RAND_360 = {1{`RANDOM}};
  _T_257_90_0 = _RAND_360[0:0];
  _RAND_361 = {1{`RANDOM}};
  _T_257_90_1 = _RAND_361[0:0];
  _RAND_362 = {1{`RANDOM}};
  _T_257_90_2 = _RAND_362[0:0];
  _RAND_363 = {1{`RANDOM}};
  _T_257_90_3 = _RAND_363[0:0];
  _RAND_364 = {1{`RANDOM}};
  _T_257_91_0 = _RAND_364[0:0];
  _RAND_365 = {1{`RANDOM}};
  _T_257_91_1 = _RAND_365[0:0];
  _RAND_366 = {1{`RANDOM}};
  _T_257_91_2 = _RAND_366[0:0];
  _RAND_367 = {1{`RANDOM}};
  _T_257_91_3 = _RAND_367[0:0];
  _RAND_368 = {1{`RANDOM}};
  _T_257_92_0 = _RAND_368[0:0];
  _RAND_369 = {1{`RANDOM}};
  _T_257_92_1 = _RAND_369[0:0];
  _RAND_370 = {1{`RANDOM}};
  _T_257_92_2 = _RAND_370[0:0];
  _RAND_371 = {1{`RANDOM}};
  _T_257_92_3 = _RAND_371[0:0];
  _RAND_372 = {1{`RANDOM}};
  _T_257_93_0 = _RAND_372[0:0];
  _RAND_373 = {1{`RANDOM}};
  _T_257_93_1 = _RAND_373[0:0];
  _RAND_374 = {1{`RANDOM}};
  _T_257_93_2 = _RAND_374[0:0];
  _RAND_375 = {1{`RANDOM}};
  _T_257_93_3 = _RAND_375[0:0];
  _RAND_376 = {1{`RANDOM}};
  _T_257_94_0 = _RAND_376[0:0];
  _RAND_377 = {1{`RANDOM}};
  _T_257_94_1 = _RAND_377[0:0];
  _RAND_378 = {1{`RANDOM}};
  _T_257_94_2 = _RAND_378[0:0];
  _RAND_379 = {1{`RANDOM}};
  _T_257_94_3 = _RAND_379[0:0];
  _RAND_380 = {1{`RANDOM}};
  _T_257_95_0 = _RAND_380[0:0];
  _RAND_381 = {1{`RANDOM}};
  _T_257_95_1 = _RAND_381[0:0];
  _RAND_382 = {1{`RANDOM}};
  _T_257_95_2 = _RAND_382[0:0];
  _RAND_383 = {1{`RANDOM}};
  _T_257_95_3 = _RAND_383[0:0];
  _RAND_384 = {1{`RANDOM}};
  _T_257_96_0 = _RAND_384[0:0];
  _RAND_385 = {1{`RANDOM}};
  _T_257_96_1 = _RAND_385[0:0];
  _RAND_386 = {1{`RANDOM}};
  _T_257_96_2 = _RAND_386[0:0];
  _RAND_387 = {1{`RANDOM}};
  _T_257_96_3 = _RAND_387[0:0];
  _RAND_388 = {1{`RANDOM}};
  _T_257_97_0 = _RAND_388[0:0];
  _RAND_389 = {1{`RANDOM}};
  _T_257_97_1 = _RAND_389[0:0];
  _RAND_390 = {1{`RANDOM}};
  _T_257_97_2 = _RAND_390[0:0];
  _RAND_391 = {1{`RANDOM}};
  _T_257_97_3 = _RAND_391[0:0];
  _RAND_392 = {1{`RANDOM}};
  _T_257_98_0 = _RAND_392[0:0];
  _RAND_393 = {1{`RANDOM}};
  _T_257_98_1 = _RAND_393[0:0];
  _RAND_394 = {1{`RANDOM}};
  _T_257_98_2 = _RAND_394[0:0];
  _RAND_395 = {1{`RANDOM}};
  _T_257_98_3 = _RAND_395[0:0];
  _RAND_396 = {1{`RANDOM}};
  _T_257_99_0 = _RAND_396[0:0];
  _RAND_397 = {1{`RANDOM}};
  _T_257_99_1 = _RAND_397[0:0];
  _RAND_398 = {1{`RANDOM}};
  _T_257_99_2 = _RAND_398[0:0];
  _RAND_399 = {1{`RANDOM}};
  _T_257_99_3 = _RAND_399[0:0];
  _RAND_400 = {1{`RANDOM}};
  _T_257_100_0 = _RAND_400[0:0];
  _RAND_401 = {1{`RANDOM}};
  _T_257_100_1 = _RAND_401[0:0];
  _RAND_402 = {1{`RANDOM}};
  _T_257_100_2 = _RAND_402[0:0];
  _RAND_403 = {1{`RANDOM}};
  _T_257_100_3 = _RAND_403[0:0];
  _RAND_404 = {1{`RANDOM}};
  _T_257_101_0 = _RAND_404[0:0];
  _RAND_405 = {1{`RANDOM}};
  _T_257_101_1 = _RAND_405[0:0];
  _RAND_406 = {1{`RANDOM}};
  _T_257_101_2 = _RAND_406[0:0];
  _RAND_407 = {1{`RANDOM}};
  _T_257_101_3 = _RAND_407[0:0];
  _RAND_408 = {1{`RANDOM}};
  _T_257_102_0 = _RAND_408[0:0];
  _RAND_409 = {1{`RANDOM}};
  _T_257_102_1 = _RAND_409[0:0];
  _RAND_410 = {1{`RANDOM}};
  _T_257_102_2 = _RAND_410[0:0];
  _RAND_411 = {1{`RANDOM}};
  _T_257_102_3 = _RAND_411[0:0];
  _RAND_412 = {1{`RANDOM}};
  _T_257_103_0 = _RAND_412[0:0];
  _RAND_413 = {1{`RANDOM}};
  _T_257_103_1 = _RAND_413[0:0];
  _RAND_414 = {1{`RANDOM}};
  _T_257_103_2 = _RAND_414[0:0];
  _RAND_415 = {1{`RANDOM}};
  _T_257_103_3 = _RAND_415[0:0];
  _RAND_416 = {1{`RANDOM}};
  _T_257_104_0 = _RAND_416[0:0];
  _RAND_417 = {1{`RANDOM}};
  _T_257_104_1 = _RAND_417[0:0];
  _RAND_418 = {1{`RANDOM}};
  _T_257_104_2 = _RAND_418[0:0];
  _RAND_419 = {1{`RANDOM}};
  _T_257_104_3 = _RAND_419[0:0];
  _RAND_420 = {1{`RANDOM}};
  _T_257_105_0 = _RAND_420[0:0];
  _RAND_421 = {1{`RANDOM}};
  _T_257_105_1 = _RAND_421[0:0];
  _RAND_422 = {1{`RANDOM}};
  _T_257_105_2 = _RAND_422[0:0];
  _RAND_423 = {1{`RANDOM}};
  _T_257_105_3 = _RAND_423[0:0];
  _RAND_424 = {1{`RANDOM}};
  _T_257_106_0 = _RAND_424[0:0];
  _RAND_425 = {1{`RANDOM}};
  _T_257_106_1 = _RAND_425[0:0];
  _RAND_426 = {1{`RANDOM}};
  _T_257_106_2 = _RAND_426[0:0];
  _RAND_427 = {1{`RANDOM}};
  _T_257_106_3 = _RAND_427[0:0];
  _RAND_428 = {1{`RANDOM}};
  _T_257_107_0 = _RAND_428[0:0];
  _RAND_429 = {1{`RANDOM}};
  _T_257_107_1 = _RAND_429[0:0];
  _RAND_430 = {1{`RANDOM}};
  _T_257_107_2 = _RAND_430[0:0];
  _RAND_431 = {1{`RANDOM}};
  _T_257_107_3 = _RAND_431[0:0];
  _RAND_432 = {1{`RANDOM}};
  _T_257_108_0 = _RAND_432[0:0];
  _RAND_433 = {1{`RANDOM}};
  _T_257_108_1 = _RAND_433[0:0];
  _RAND_434 = {1{`RANDOM}};
  _T_257_108_2 = _RAND_434[0:0];
  _RAND_435 = {1{`RANDOM}};
  _T_257_108_3 = _RAND_435[0:0];
  _RAND_436 = {1{`RANDOM}};
  _T_257_109_0 = _RAND_436[0:0];
  _RAND_437 = {1{`RANDOM}};
  _T_257_109_1 = _RAND_437[0:0];
  _RAND_438 = {1{`RANDOM}};
  _T_257_109_2 = _RAND_438[0:0];
  _RAND_439 = {1{`RANDOM}};
  _T_257_109_3 = _RAND_439[0:0];
  _RAND_440 = {1{`RANDOM}};
  _T_257_110_0 = _RAND_440[0:0];
  _RAND_441 = {1{`RANDOM}};
  _T_257_110_1 = _RAND_441[0:0];
  _RAND_442 = {1{`RANDOM}};
  _T_257_110_2 = _RAND_442[0:0];
  _RAND_443 = {1{`RANDOM}};
  _T_257_110_3 = _RAND_443[0:0];
  _RAND_444 = {1{`RANDOM}};
  _T_257_111_0 = _RAND_444[0:0];
  _RAND_445 = {1{`RANDOM}};
  _T_257_111_1 = _RAND_445[0:0];
  _RAND_446 = {1{`RANDOM}};
  _T_257_111_2 = _RAND_446[0:0];
  _RAND_447 = {1{`RANDOM}};
  _T_257_111_3 = _RAND_447[0:0];
  _RAND_448 = {1{`RANDOM}};
  _T_257_112_0 = _RAND_448[0:0];
  _RAND_449 = {1{`RANDOM}};
  _T_257_112_1 = _RAND_449[0:0];
  _RAND_450 = {1{`RANDOM}};
  _T_257_112_2 = _RAND_450[0:0];
  _RAND_451 = {1{`RANDOM}};
  _T_257_112_3 = _RAND_451[0:0];
  _RAND_452 = {1{`RANDOM}};
  _T_257_113_0 = _RAND_452[0:0];
  _RAND_453 = {1{`RANDOM}};
  _T_257_113_1 = _RAND_453[0:0];
  _RAND_454 = {1{`RANDOM}};
  _T_257_113_2 = _RAND_454[0:0];
  _RAND_455 = {1{`RANDOM}};
  _T_257_113_3 = _RAND_455[0:0];
  _RAND_456 = {1{`RANDOM}};
  _T_257_114_0 = _RAND_456[0:0];
  _RAND_457 = {1{`RANDOM}};
  _T_257_114_1 = _RAND_457[0:0];
  _RAND_458 = {1{`RANDOM}};
  _T_257_114_2 = _RAND_458[0:0];
  _RAND_459 = {1{`RANDOM}};
  _T_257_114_3 = _RAND_459[0:0];
  _RAND_460 = {1{`RANDOM}};
  _T_257_115_0 = _RAND_460[0:0];
  _RAND_461 = {1{`RANDOM}};
  _T_257_115_1 = _RAND_461[0:0];
  _RAND_462 = {1{`RANDOM}};
  _T_257_115_2 = _RAND_462[0:0];
  _RAND_463 = {1{`RANDOM}};
  _T_257_115_3 = _RAND_463[0:0];
  _RAND_464 = {1{`RANDOM}};
  _T_257_116_0 = _RAND_464[0:0];
  _RAND_465 = {1{`RANDOM}};
  _T_257_116_1 = _RAND_465[0:0];
  _RAND_466 = {1{`RANDOM}};
  _T_257_116_2 = _RAND_466[0:0];
  _RAND_467 = {1{`RANDOM}};
  _T_257_116_3 = _RAND_467[0:0];
  _RAND_468 = {1{`RANDOM}};
  _T_257_117_0 = _RAND_468[0:0];
  _RAND_469 = {1{`RANDOM}};
  _T_257_117_1 = _RAND_469[0:0];
  _RAND_470 = {1{`RANDOM}};
  _T_257_117_2 = _RAND_470[0:0];
  _RAND_471 = {1{`RANDOM}};
  _T_257_117_3 = _RAND_471[0:0];
  _RAND_472 = {1{`RANDOM}};
  _T_257_118_0 = _RAND_472[0:0];
  _RAND_473 = {1{`RANDOM}};
  _T_257_118_1 = _RAND_473[0:0];
  _RAND_474 = {1{`RANDOM}};
  _T_257_118_2 = _RAND_474[0:0];
  _RAND_475 = {1{`RANDOM}};
  _T_257_118_3 = _RAND_475[0:0];
  _RAND_476 = {1{`RANDOM}};
  _T_257_119_0 = _RAND_476[0:0];
  _RAND_477 = {1{`RANDOM}};
  _T_257_119_1 = _RAND_477[0:0];
  _RAND_478 = {1{`RANDOM}};
  _T_257_119_2 = _RAND_478[0:0];
  _RAND_479 = {1{`RANDOM}};
  _T_257_119_3 = _RAND_479[0:0];
  _RAND_480 = {1{`RANDOM}};
  _T_257_120_0 = _RAND_480[0:0];
  _RAND_481 = {1{`RANDOM}};
  _T_257_120_1 = _RAND_481[0:0];
  _RAND_482 = {1{`RANDOM}};
  _T_257_120_2 = _RAND_482[0:0];
  _RAND_483 = {1{`RANDOM}};
  _T_257_120_3 = _RAND_483[0:0];
  _RAND_484 = {1{`RANDOM}};
  _T_257_121_0 = _RAND_484[0:0];
  _RAND_485 = {1{`RANDOM}};
  _T_257_121_1 = _RAND_485[0:0];
  _RAND_486 = {1{`RANDOM}};
  _T_257_121_2 = _RAND_486[0:0];
  _RAND_487 = {1{`RANDOM}};
  _T_257_121_3 = _RAND_487[0:0];
  _RAND_488 = {1{`RANDOM}};
  _T_257_122_0 = _RAND_488[0:0];
  _RAND_489 = {1{`RANDOM}};
  _T_257_122_1 = _RAND_489[0:0];
  _RAND_490 = {1{`RANDOM}};
  _T_257_122_2 = _RAND_490[0:0];
  _RAND_491 = {1{`RANDOM}};
  _T_257_122_3 = _RAND_491[0:0];
  _RAND_492 = {1{`RANDOM}};
  _T_257_123_0 = _RAND_492[0:0];
  _RAND_493 = {1{`RANDOM}};
  _T_257_123_1 = _RAND_493[0:0];
  _RAND_494 = {1{`RANDOM}};
  _T_257_123_2 = _RAND_494[0:0];
  _RAND_495 = {1{`RANDOM}};
  _T_257_123_3 = _RAND_495[0:0];
  _RAND_496 = {1{`RANDOM}};
  _T_257_124_0 = _RAND_496[0:0];
  _RAND_497 = {1{`RANDOM}};
  _T_257_124_1 = _RAND_497[0:0];
  _RAND_498 = {1{`RANDOM}};
  _T_257_124_2 = _RAND_498[0:0];
  _RAND_499 = {1{`RANDOM}};
  _T_257_124_3 = _RAND_499[0:0];
  _RAND_500 = {1{`RANDOM}};
  _T_257_125_0 = _RAND_500[0:0];
  _RAND_501 = {1{`RANDOM}};
  _T_257_125_1 = _RAND_501[0:0];
  _RAND_502 = {1{`RANDOM}};
  _T_257_125_2 = _RAND_502[0:0];
  _RAND_503 = {1{`RANDOM}};
  _T_257_125_3 = _RAND_503[0:0];
  _RAND_504 = {1{`RANDOM}};
  _T_257_126_0 = _RAND_504[0:0];
  _RAND_505 = {1{`RANDOM}};
  _T_257_126_1 = _RAND_505[0:0];
  _RAND_506 = {1{`RANDOM}};
  _T_257_126_2 = _RAND_506[0:0];
  _RAND_507 = {1{`RANDOM}};
  _T_257_126_3 = _RAND_507[0:0];
  _RAND_508 = {1{`RANDOM}};
  _T_257_127_0 = _RAND_508[0:0];
  _RAND_509 = {1{`RANDOM}};
  _T_257_127_1 = _RAND_509[0:0];
  _RAND_510 = {1{`RANDOM}};
  _T_257_127_2 = _RAND_510[0:0];
  _RAND_511 = {1{`RANDOM}};
  _T_257_127_3 = _RAND_511[0:0];
  _RAND_512 = {1{`RANDOM}};
  _T_257_128_0 = _RAND_512[0:0];
  _RAND_513 = {1{`RANDOM}};
  _T_257_128_1 = _RAND_513[0:0];
  _RAND_514 = {1{`RANDOM}};
  _T_257_128_2 = _RAND_514[0:0];
  _RAND_515 = {1{`RANDOM}};
  _T_257_128_3 = _RAND_515[0:0];
  _RAND_516 = {1{`RANDOM}};
  _T_257_129_0 = _RAND_516[0:0];
  _RAND_517 = {1{`RANDOM}};
  _T_257_129_1 = _RAND_517[0:0];
  _RAND_518 = {1{`RANDOM}};
  _T_257_129_2 = _RAND_518[0:0];
  _RAND_519 = {1{`RANDOM}};
  _T_257_129_3 = _RAND_519[0:0];
  _RAND_520 = {1{`RANDOM}};
  _T_257_130_0 = _RAND_520[0:0];
  _RAND_521 = {1{`RANDOM}};
  _T_257_130_1 = _RAND_521[0:0];
  _RAND_522 = {1{`RANDOM}};
  _T_257_130_2 = _RAND_522[0:0];
  _RAND_523 = {1{`RANDOM}};
  _T_257_130_3 = _RAND_523[0:0];
  _RAND_524 = {1{`RANDOM}};
  _T_257_131_0 = _RAND_524[0:0];
  _RAND_525 = {1{`RANDOM}};
  _T_257_131_1 = _RAND_525[0:0];
  _RAND_526 = {1{`RANDOM}};
  _T_257_131_2 = _RAND_526[0:0];
  _RAND_527 = {1{`RANDOM}};
  _T_257_131_3 = _RAND_527[0:0];
  _RAND_528 = {1{`RANDOM}};
  _T_257_132_0 = _RAND_528[0:0];
  _RAND_529 = {1{`RANDOM}};
  _T_257_132_1 = _RAND_529[0:0];
  _RAND_530 = {1{`RANDOM}};
  _T_257_132_2 = _RAND_530[0:0];
  _RAND_531 = {1{`RANDOM}};
  _T_257_132_3 = _RAND_531[0:0];
  _RAND_532 = {1{`RANDOM}};
  _T_257_133_0 = _RAND_532[0:0];
  _RAND_533 = {1{`RANDOM}};
  _T_257_133_1 = _RAND_533[0:0];
  _RAND_534 = {1{`RANDOM}};
  _T_257_133_2 = _RAND_534[0:0];
  _RAND_535 = {1{`RANDOM}};
  _T_257_133_3 = _RAND_535[0:0];
  _RAND_536 = {1{`RANDOM}};
  _T_257_134_0 = _RAND_536[0:0];
  _RAND_537 = {1{`RANDOM}};
  _T_257_134_1 = _RAND_537[0:0];
  _RAND_538 = {1{`RANDOM}};
  _T_257_134_2 = _RAND_538[0:0];
  _RAND_539 = {1{`RANDOM}};
  _T_257_134_3 = _RAND_539[0:0];
  _RAND_540 = {1{`RANDOM}};
  _T_257_135_0 = _RAND_540[0:0];
  _RAND_541 = {1{`RANDOM}};
  _T_257_135_1 = _RAND_541[0:0];
  _RAND_542 = {1{`RANDOM}};
  _T_257_135_2 = _RAND_542[0:0];
  _RAND_543 = {1{`RANDOM}};
  _T_257_135_3 = _RAND_543[0:0];
  _RAND_544 = {1{`RANDOM}};
  _T_257_136_0 = _RAND_544[0:0];
  _RAND_545 = {1{`RANDOM}};
  _T_257_136_1 = _RAND_545[0:0];
  _RAND_546 = {1{`RANDOM}};
  _T_257_136_2 = _RAND_546[0:0];
  _RAND_547 = {1{`RANDOM}};
  _T_257_136_3 = _RAND_547[0:0];
  _RAND_548 = {1{`RANDOM}};
  _T_257_137_0 = _RAND_548[0:0];
  _RAND_549 = {1{`RANDOM}};
  _T_257_137_1 = _RAND_549[0:0];
  _RAND_550 = {1{`RANDOM}};
  _T_257_137_2 = _RAND_550[0:0];
  _RAND_551 = {1{`RANDOM}};
  _T_257_137_3 = _RAND_551[0:0];
  _RAND_552 = {1{`RANDOM}};
  _T_257_138_0 = _RAND_552[0:0];
  _RAND_553 = {1{`RANDOM}};
  _T_257_138_1 = _RAND_553[0:0];
  _RAND_554 = {1{`RANDOM}};
  _T_257_138_2 = _RAND_554[0:0];
  _RAND_555 = {1{`RANDOM}};
  _T_257_138_3 = _RAND_555[0:0];
  _RAND_556 = {1{`RANDOM}};
  _T_257_139_0 = _RAND_556[0:0];
  _RAND_557 = {1{`RANDOM}};
  _T_257_139_1 = _RAND_557[0:0];
  _RAND_558 = {1{`RANDOM}};
  _T_257_139_2 = _RAND_558[0:0];
  _RAND_559 = {1{`RANDOM}};
  _T_257_139_3 = _RAND_559[0:0];
  _RAND_560 = {1{`RANDOM}};
  _T_257_140_0 = _RAND_560[0:0];
  _RAND_561 = {1{`RANDOM}};
  _T_257_140_1 = _RAND_561[0:0];
  _RAND_562 = {1{`RANDOM}};
  _T_257_140_2 = _RAND_562[0:0];
  _RAND_563 = {1{`RANDOM}};
  _T_257_140_3 = _RAND_563[0:0];
  _RAND_564 = {1{`RANDOM}};
  _T_257_141_0 = _RAND_564[0:0];
  _RAND_565 = {1{`RANDOM}};
  _T_257_141_1 = _RAND_565[0:0];
  _RAND_566 = {1{`RANDOM}};
  _T_257_141_2 = _RAND_566[0:0];
  _RAND_567 = {1{`RANDOM}};
  _T_257_141_3 = _RAND_567[0:0];
  _RAND_568 = {1{`RANDOM}};
  _T_257_142_0 = _RAND_568[0:0];
  _RAND_569 = {1{`RANDOM}};
  _T_257_142_1 = _RAND_569[0:0];
  _RAND_570 = {1{`RANDOM}};
  _T_257_142_2 = _RAND_570[0:0];
  _RAND_571 = {1{`RANDOM}};
  _T_257_142_3 = _RAND_571[0:0];
  _RAND_572 = {1{`RANDOM}};
  _T_257_143_0 = _RAND_572[0:0];
  _RAND_573 = {1{`RANDOM}};
  _T_257_143_1 = _RAND_573[0:0];
  _RAND_574 = {1{`RANDOM}};
  _T_257_143_2 = _RAND_574[0:0];
  _RAND_575 = {1{`RANDOM}};
  _T_257_143_3 = _RAND_575[0:0];
  _RAND_576 = {1{`RANDOM}};
  _T_257_144_0 = _RAND_576[0:0];
  _RAND_577 = {1{`RANDOM}};
  _T_257_144_1 = _RAND_577[0:0];
  _RAND_578 = {1{`RANDOM}};
  _T_257_144_2 = _RAND_578[0:0];
  _RAND_579 = {1{`RANDOM}};
  _T_257_144_3 = _RAND_579[0:0];
  _RAND_580 = {1{`RANDOM}};
  _T_257_145_0 = _RAND_580[0:0];
  _RAND_581 = {1{`RANDOM}};
  _T_257_145_1 = _RAND_581[0:0];
  _RAND_582 = {1{`RANDOM}};
  _T_257_145_2 = _RAND_582[0:0];
  _RAND_583 = {1{`RANDOM}};
  _T_257_145_3 = _RAND_583[0:0];
  _RAND_584 = {1{`RANDOM}};
  _T_257_146_0 = _RAND_584[0:0];
  _RAND_585 = {1{`RANDOM}};
  _T_257_146_1 = _RAND_585[0:0];
  _RAND_586 = {1{`RANDOM}};
  _T_257_146_2 = _RAND_586[0:0];
  _RAND_587 = {1{`RANDOM}};
  _T_257_146_3 = _RAND_587[0:0];
  _RAND_588 = {1{`RANDOM}};
  _T_257_147_0 = _RAND_588[0:0];
  _RAND_589 = {1{`RANDOM}};
  _T_257_147_1 = _RAND_589[0:0];
  _RAND_590 = {1{`RANDOM}};
  _T_257_147_2 = _RAND_590[0:0];
  _RAND_591 = {1{`RANDOM}};
  _T_257_147_3 = _RAND_591[0:0];
  _RAND_592 = {1{`RANDOM}};
  _T_257_148_0 = _RAND_592[0:0];
  _RAND_593 = {1{`RANDOM}};
  _T_257_148_1 = _RAND_593[0:0];
  _RAND_594 = {1{`RANDOM}};
  _T_257_148_2 = _RAND_594[0:0];
  _RAND_595 = {1{`RANDOM}};
  _T_257_148_3 = _RAND_595[0:0];
  _RAND_596 = {1{`RANDOM}};
  _T_257_149_0 = _RAND_596[0:0];
  _RAND_597 = {1{`RANDOM}};
  _T_257_149_1 = _RAND_597[0:0];
  _RAND_598 = {1{`RANDOM}};
  _T_257_149_2 = _RAND_598[0:0];
  _RAND_599 = {1{`RANDOM}};
  _T_257_149_3 = _RAND_599[0:0];
  _RAND_600 = {1{`RANDOM}};
  _T_257_150_0 = _RAND_600[0:0];
  _RAND_601 = {1{`RANDOM}};
  _T_257_150_1 = _RAND_601[0:0];
  _RAND_602 = {1{`RANDOM}};
  _T_257_150_2 = _RAND_602[0:0];
  _RAND_603 = {1{`RANDOM}};
  _T_257_150_3 = _RAND_603[0:0];
  _RAND_604 = {1{`RANDOM}};
  _T_257_151_0 = _RAND_604[0:0];
  _RAND_605 = {1{`RANDOM}};
  _T_257_151_1 = _RAND_605[0:0];
  _RAND_606 = {1{`RANDOM}};
  _T_257_151_2 = _RAND_606[0:0];
  _RAND_607 = {1{`RANDOM}};
  _T_257_151_3 = _RAND_607[0:0];
  _RAND_608 = {1{`RANDOM}};
  _T_257_152_0 = _RAND_608[0:0];
  _RAND_609 = {1{`RANDOM}};
  _T_257_152_1 = _RAND_609[0:0];
  _RAND_610 = {1{`RANDOM}};
  _T_257_152_2 = _RAND_610[0:0];
  _RAND_611 = {1{`RANDOM}};
  _T_257_152_3 = _RAND_611[0:0];
  _RAND_612 = {1{`RANDOM}};
  _T_257_153_0 = _RAND_612[0:0];
  _RAND_613 = {1{`RANDOM}};
  _T_257_153_1 = _RAND_613[0:0];
  _RAND_614 = {1{`RANDOM}};
  _T_257_153_2 = _RAND_614[0:0];
  _RAND_615 = {1{`RANDOM}};
  _T_257_153_3 = _RAND_615[0:0];
  _RAND_616 = {1{`RANDOM}};
  _T_257_154_0 = _RAND_616[0:0];
  _RAND_617 = {1{`RANDOM}};
  _T_257_154_1 = _RAND_617[0:0];
  _RAND_618 = {1{`RANDOM}};
  _T_257_154_2 = _RAND_618[0:0];
  _RAND_619 = {1{`RANDOM}};
  _T_257_154_3 = _RAND_619[0:0];
  _RAND_620 = {1{`RANDOM}};
  _T_257_155_0 = _RAND_620[0:0];
  _RAND_621 = {1{`RANDOM}};
  _T_257_155_1 = _RAND_621[0:0];
  _RAND_622 = {1{`RANDOM}};
  _T_257_155_2 = _RAND_622[0:0];
  _RAND_623 = {1{`RANDOM}};
  _T_257_155_3 = _RAND_623[0:0];
  _RAND_624 = {1{`RANDOM}};
  _T_257_156_0 = _RAND_624[0:0];
  _RAND_625 = {1{`RANDOM}};
  _T_257_156_1 = _RAND_625[0:0];
  _RAND_626 = {1{`RANDOM}};
  _T_257_156_2 = _RAND_626[0:0];
  _RAND_627 = {1{`RANDOM}};
  _T_257_156_3 = _RAND_627[0:0];
  _RAND_628 = {1{`RANDOM}};
  _T_257_157_0 = _RAND_628[0:0];
  _RAND_629 = {1{`RANDOM}};
  _T_257_157_1 = _RAND_629[0:0];
  _RAND_630 = {1{`RANDOM}};
  _T_257_157_2 = _RAND_630[0:0];
  _RAND_631 = {1{`RANDOM}};
  _T_257_157_3 = _RAND_631[0:0];
  _RAND_632 = {1{`RANDOM}};
  _T_257_158_0 = _RAND_632[0:0];
  _RAND_633 = {1{`RANDOM}};
  _T_257_158_1 = _RAND_633[0:0];
  _RAND_634 = {1{`RANDOM}};
  _T_257_158_2 = _RAND_634[0:0];
  _RAND_635 = {1{`RANDOM}};
  _T_257_158_3 = _RAND_635[0:0];
  _RAND_636 = {1{`RANDOM}};
  _T_257_159_0 = _RAND_636[0:0];
  _RAND_637 = {1{`RANDOM}};
  _T_257_159_1 = _RAND_637[0:0];
  _RAND_638 = {1{`RANDOM}};
  _T_257_159_2 = _RAND_638[0:0];
  _RAND_639 = {1{`RANDOM}};
  _T_257_159_3 = _RAND_639[0:0];
  _RAND_640 = {1{`RANDOM}};
  _T_257_160_0 = _RAND_640[0:0];
  _RAND_641 = {1{`RANDOM}};
  _T_257_160_1 = _RAND_641[0:0];
  _RAND_642 = {1{`RANDOM}};
  _T_257_160_2 = _RAND_642[0:0];
  _RAND_643 = {1{`RANDOM}};
  _T_257_160_3 = _RAND_643[0:0];
  _RAND_644 = {1{`RANDOM}};
  _T_257_161_0 = _RAND_644[0:0];
  _RAND_645 = {1{`RANDOM}};
  _T_257_161_1 = _RAND_645[0:0];
  _RAND_646 = {1{`RANDOM}};
  _T_257_161_2 = _RAND_646[0:0];
  _RAND_647 = {1{`RANDOM}};
  _T_257_161_3 = _RAND_647[0:0];
  _RAND_648 = {1{`RANDOM}};
  _T_257_162_0 = _RAND_648[0:0];
  _RAND_649 = {1{`RANDOM}};
  _T_257_162_1 = _RAND_649[0:0];
  _RAND_650 = {1{`RANDOM}};
  _T_257_162_2 = _RAND_650[0:0];
  _RAND_651 = {1{`RANDOM}};
  _T_257_162_3 = _RAND_651[0:0];
  _RAND_652 = {1{`RANDOM}};
  _T_257_163_0 = _RAND_652[0:0];
  _RAND_653 = {1{`RANDOM}};
  _T_257_163_1 = _RAND_653[0:0];
  _RAND_654 = {1{`RANDOM}};
  _T_257_163_2 = _RAND_654[0:0];
  _RAND_655 = {1{`RANDOM}};
  _T_257_163_3 = _RAND_655[0:0];
  _RAND_656 = {1{`RANDOM}};
  _T_257_164_0 = _RAND_656[0:0];
  _RAND_657 = {1{`RANDOM}};
  _T_257_164_1 = _RAND_657[0:0];
  _RAND_658 = {1{`RANDOM}};
  _T_257_164_2 = _RAND_658[0:0];
  _RAND_659 = {1{`RANDOM}};
  _T_257_164_3 = _RAND_659[0:0];
  _RAND_660 = {1{`RANDOM}};
  _T_257_165_0 = _RAND_660[0:0];
  _RAND_661 = {1{`RANDOM}};
  _T_257_165_1 = _RAND_661[0:0];
  _RAND_662 = {1{`RANDOM}};
  _T_257_165_2 = _RAND_662[0:0];
  _RAND_663 = {1{`RANDOM}};
  _T_257_165_3 = _RAND_663[0:0];
  _RAND_664 = {1{`RANDOM}};
  _T_257_166_0 = _RAND_664[0:0];
  _RAND_665 = {1{`RANDOM}};
  _T_257_166_1 = _RAND_665[0:0];
  _RAND_666 = {1{`RANDOM}};
  _T_257_166_2 = _RAND_666[0:0];
  _RAND_667 = {1{`RANDOM}};
  _T_257_166_3 = _RAND_667[0:0];
  _RAND_668 = {1{`RANDOM}};
  _T_257_167_0 = _RAND_668[0:0];
  _RAND_669 = {1{`RANDOM}};
  _T_257_167_1 = _RAND_669[0:0];
  _RAND_670 = {1{`RANDOM}};
  _T_257_167_2 = _RAND_670[0:0];
  _RAND_671 = {1{`RANDOM}};
  _T_257_167_3 = _RAND_671[0:0];
  _RAND_672 = {1{`RANDOM}};
  _T_257_168_0 = _RAND_672[0:0];
  _RAND_673 = {1{`RANDOM}};
  _T_257_168_1 = _RAND_673[0:0];
  _RAND_674 = {1{`RANDOM}};
  _T_257_168_2 = _RAND_674[0:0];
  _RAND_675 = {1{`RANDOM}};
  _T_257_168_3 = _RAND_675[0:0];
  _RAND_676 = {1{`RANDOM}};
  _T_257_169_0 = _RAND_676[0:0];
  _RAND_677 = {1{`RANDOM}};
  _T_257_169_1 = _RAND_677[0:0];
  _RAND_678 = {1{`RANDOM}};
  _T_257_169_2 = _RAND_678[0:0];
  _RAND_679 = {1{`RANDOM}};
  _T_257_169_3 = _RAND_679[0:0];
  _RAND_680 = {1{`RANDOM}};
  _T_257_170_0 = _RAND_680[0:0];
  _RAND_681 = {1{`RANDOM}};
  _T_257_170_1 = _RAND_681[0:0];
  _RAND_682 = {1{`RANDOM}};
  _T_257_170_2 = _RAND_682[0:0];
  _RAND_683 = {1{`RANDOM}};
  _T_257_170_3 = _RAND_683[0:0];
  _RAND_684 = {1{`RANDOM}};
  _T_257_171_0 = _RAND_684[0:0];
  _RAND_685 = {1{`RANDOM}};
  _T_257_171_1 = _RAND_685[0:0];
  _RAND_686 = {1{`RANDOM}};
  _T_257_171_2 = _RAND_686[0:0];
  _RAND_687 = {1{`RANDOM}};
  _T_257_171_3 = _RAND_687[0:0];
  _RAND_688 = {1{`RANDOM}};
  _T_257_172_0 = _RAND_688[0:0];
  _RAND_689 = {1{`RANDOM}};
  _T_257_172_1 = _RAND_689[0:0];
  _RAND_690 = {1{`RANDOM}};
  _T_257_172_2 = _RAND_690[0:0];
  _RAND_691 = {1{`RANDOM}};
  _T_257_172_3 = _RAND_691[0:0];
  _RAND_692 = {1{`RANDOM}};
  _T_257_173_0 = _RAND_692[0:0];
  _RAND_693 = {1{`RANDOM}};
  _T_257_173_1 = _RAND_693[0:0];
  _RAND_694 = {1{`RANDOM}};
  _T_257_173_2 = _RAND_694[0:0];
  _RAND_695 = {1{`RANDOM}};
  _T_257_173_3 = _RAND_695[0:0];
  _RAND_696 = {1{`RANDOM}};
  _T_257_174_0 = _RAND_696[0:0];
  _RAND_697 = {1{`RANDOM}};
  _T_257_174_1 = _RAND_697[0:0];
  _RAND_698 = {1{`RANDOM}};
  _T_257_174_2 = _RAND_698[0:0];
  _RAND_699 = {1{`RANDOM}};
  _T_257_174_3 = _RAND_699[0:0];
  _RAND_700 = {1{`RANDOM}};
  _T_257_175_0 = _RAND_700[0:0];
  _RAND_701 = {1{`RANDOM}};
  _T_257_175_1 = _RAND_701[0:0];
  _RAND_702 = {1{`RANDOM}};
  _T_257_175_2 = _RAND_702[0:0];
  _RAND_703 = {1{`RANDOM}};
  _T_257_175_3 = _RAND_703[0:0];
  _RAND_704 = {1{`RANDOM}};
  _T_257_176_0 = _RAND_704[0:0];
  _RAND_705 = {1{`RANDOM}};
  _T_257_176_1 = _RAND_705[0:0];
  _RAND_706 = {1{`RANDOM}};
  _T_257_176_2 = _RAND_706[0:0];
  _RAND_707 = {1{`RANDOM}};
  _T_257_176_3 = _RAND_707[0:0];
  _RAND_708 = {1{`RANDOM}};
  _T_257_177_0 = _RAND_708[0:0];
  _RAND_709 = {1{`RANDOM}};
  _T_257_177_1 = _RAND_709[0:0];
  _RAND_710 = {1{`RANDOM}};
  _T_257_177_2 = _RAND_710[0:0];
  _RAND_711 = {1{`RANDOM}};
  _T_257_177_3 = _RAND_711[0:0];
  _RAND_712 = {1{`RANDOM}};
  _T_257_178_0 = _RAND_712[0:0];
  _RAND_713 = {1{`RANDOM}};
  _T_257_178_1 = _RAND_713[0:0];
  _RAND_714 = {1{`RANDOM}};
  _T_257_178_2 = _RAND_714[0:0];
  _RAND_715 = {1{`RANDOM}};
  _T_257_178_3 = _RAND_715[0:0];
  _RAND_716 = {1{`RANDOM}};
  _T_257_179_0 = _RAND_716[0:0];
  _RAND_717 = {1{`RANDOM}};
  _T_257_179_1 = _RAND_717[0:0];
  _RAND_718 = {1{`RANDOM}};
  _T_257_179_2 = _RAND_718[0:0];
  _RAND_719 = {1{`RANDOM}};
  _T_257_179_3 = _RAND_719[0:0];
  _RAND_720 = {1{`RANDOM}};
  _T_257_180_0 = _RAND_720[0:0];
  _RAND_721 = {1{`RANDOM}};
  _T_257_180_1 = _RAND_721[0:0];
  _RAND_722 = {1{`RANDOM}};
  _T_257_180_2 = _RAND_722[0:0];
  _RAND_723 = {1{`RANDOM}};
  _T_257_180_3 = _RAND_723[0:0];
  _RAND_724 = {1{`RANDOM}};
  _T_257_181_0 = _RAND_724[0:0];
  _RAND_725 = {1{`RANDOM}};
  _T_257_181_1 = _RAND_725[0:0];
  _RAND_726 = {1{`RANDOM}};
  _T_257_181_2 = _RAND_726[0:0];
  _RAND_727 = {1{`RANDOM}};
  _T_257_181_3 = _RAND_727[0:0];
  _RAND_728 = {1{`RANDOM}};
  _T_257_182_0 = _RAND_728[0:0];
  _RAND_729 = {1{`RANDOM}};
  _T_257_182_1 = _RAND_729[0:0];
  _RAND_730 = {1{`RANDOM}};
  _T_257_182_2 = _RAND_730[0:0];
  _RAND_731 = {1{`RANDOM}};
  _T_257_182_3 = _RAND_731[0:0];
  _RAND_732 = {1{`RANDOM}};
  _T_257_183_0 = _RAND_732[0:0];
  _RAND_733 = {1{`RANDOM}};
  _T_257_183_1 = _RAND_733[0:0];
  _RAND_734 = {1{`RANDOM}};
  _T_257_183_2 = _RAND_734[0:0];
  _RAND_735 = {1{`RANDOM}};
  _T_257_183_3 = _RAND_735[0:0];
  _RAND_736 = {1{`RANDOM}};
  _T_257_184_0 = _RAND_736[0:0];
  _RAND_737 = {1{`RANDOM}};
  _T_257_184_1 = _RAND_737[0:0];
  _RAND_738 = {1{`RANDOM}};
  _T_257_184_2 = _RAND_738[0:0];
  _RAND_739 = {1{`RANDOM}};
  _T_257_184_3 = _RAND_739[0:0];
  _RAND_740 = {1{`RANDOM}};
  _T_257_185_0 = _RAND_740[0:0];
  _RAND_741 = {1{`RANDOM}};
  _T_257_185_1 = _RAND_741[0:0];
  _RAND_742 = {1{`RANDOM}};
  _T_257_185_2 = _RAND_742[0:0];
  _RAND_743 = {1{`RANDOM}};
  _T_257_185_3 = _RAND_743[0:0];
  _RAND_744 = {1{`RANDOM}};
  _T_257_186_0 = _RAND_744[0:0];
  _RAND_745 = {1{`RANDOM}};
  _T_257_186_1 = _RAND_745[0:0];
  _RAND_746 = {1{`RANDOM}};
  _T_257_186_2 = _RAND_746[0:0];
  _RAND_747 = {1{`RANDOM}};
  _T_257_186_3 = _RAND_747[0:0];
  _RAND_748 = {1{`RANDOM}};
  _T_257_187_0 = _RAND_748[0:0];
  _RAND_749 = {1{`RANDOM}};
  _T_257_187_1 = _RAND_749[0:0];
  _RAND_750 = {1{`RANDOM}};
  _T_257_187_2 = _RAND_750[0:0];
  _RAND_751 = {1{`RANDOM}};
  _T_257_187_3 = _RAND_751[0:0];
  _RAND_752 = {1{`RANDOM}};
  _T_257_188_0 = _RAND_752[0:0];
  _RAND_753 = {1{`RANDOM}};
  _T_257_188_1 = _RAND_753[0:0];
  _RAND_754 = {1{`RANDOM}};
  _T_257_188_2 = _RAND_754[0:0];
  _RAND_755 = {1{`RANDOM}};
  _T_257_188_3 = _RAND_755[0:0];
  _RAND_756 = {1{`RANDOM}};
  _T_257_189_0 = _RAND_756[0:0];
  _RAND_757 = {1{`RANDOM}};
  _T_257_189_1 = _RAND_757[0:0];
  _RAND_758 = {1{`RANDOM}};
  _T_257_189_2 = _RAND_758[0:0];
  _RAND_759 = {1{`RANDOM}};
  _T_257_189_3 = _RAND_759[0:0];
  _RAND_760 = {1{`RANDOM}};
  _T_257_190_0 = _RAND_760[0:0];
  _RAND_761 = {1{`RANDOM}};
  _T_257_190_1 = _RAND_761[0:0];
  _RAND_762 = {1{`RANDOM}};
  _T_257_190_2 = _RAND_762[0:0];
  _RAND_763 = {1{`RANDOM}};
  _T_257_190_3 = _RAND_763[0:0];
  _RAND_764 = {1{`RANDOM}};
  _T_257_191_0 = _RAND_764[0:0];
  _RAND_765 = {1{`RANDOM}};
  _T_257_191_1 = _RAND_765[0:0];
  _RAND_766 = {1{`RANDOM}};
  _T_257_191_2 = _RAND_766[0:0];
  _RAND_767 = {1{`RANDOM}};
  _T_257_191_3 = _RAND_767[0:0];
  _RAND_768 = {1{`RANDOM}};
  _T_257_192_0 = _RAND_768[0:0];
  _RAND_769 = {1{`RANDOM}};
  _T_257_192_1 = _RAND_769[0:0];
  _RAND_770 = {1{`RANDOM}};
  _T_257_192_2 = _RAND_770[0:0];
  _RAND_771 = {1{`RANDOM}};
  _T_257_192_3 = _RAND_771[0:0];
  _RAND_772 = {1{`RANDOM}};
  _T_257_193_0 = _RAND_772[0:0];
  _RAND_773 = {1{`RANDOM}};
  _T_257_193_1 = _RAND_773[0:0];
  _RAND_774 = {1{`RANDOM}};
  _T_257_193_2 = _RAND_774[0:0];
  _RAND_775 = {1{`RANDOM}};
  _T_257_193_3 = _RAND_775[0:0];
  _RAND_776 = {1{`RANDOM}};
  _T_257_194_0 = _RAND_776[0:0];
  _RAND_777 = {1{`RANDOM}};
  _T_257_194_1 = _RAND_777[0:0];
  _RAND_778 = {1{`RANDOM}};
  _T_257_194_2 = _RAND_778[0:0];
  _RAND_779 = {1{`RANDOM}};
  _T_257_194_3 = _RAND_779[0:0];
  _RAND_780 = {1{`RANDOM}};
  _T_257_195_0 = _RAND_780[0:0];
  _RAND_781 = {1{`RANDOM}};
  _T_257_195_1 = _RAND_781[0:0];
  _RAND_782 = {1{`RANDOM}};
  _T_257_195_2 = _RAND_782[0:0];
  _RAND_783 = {1{`RANDOM}};
  _T_257_195_3 = _RAND_783[0:0];
  _RAND_784 = {1{`RANDOM}};
  _T_257_196_0 = _RAND_784[0:0];
  _RAND_785 = {1{`RANDOM}};
  _T_257_196_1 = _RAND_785[0:0];
  _RAND_786 = {1{`RANDOM}};
  _T_257_196_2 = _RAND_786[0:0];
  _RAND_787 = {1{`RANDOM}};
  _T_257_196_3 = _RAND_787[0:0];
  _RAND_788 = {1{`RANDOM}};
  _T_257_197_0 = _RAND_788[0:0];
  _RAND_789 = {1{`RANDOM}};
  _T_257_197_1 = _RAND_789[0:0];
  _RAND_790 = {1{`RANDOM}};
  _T_257_197_2 = _RAND_790[0:0];
  _RAND_791 = {1{`RANDOM}};
  _T_257_197_3 = _RAND_791[0:0];
  _RAND_792 = {1{`RANDOM}};
  _T_257_198_0 = _RAND_792[0:0];
  _RAND_793 = {1{`RANDOM}};
  _T_257_198_1 = _RAND_793[0:0];
  _RAND_794 = {1{`RANDOM}};
  _T_257_198_2 = _RAND_794[0:0];
  _RAND_795 = {1{`RANDOM}};
  _T_257_198_3 = _RAND_795[0:0];
  _RAND_796 = {1{`RANDOM}};
  _T_257_199_0 = _RAND_796[0:0];
  _RAND_797 = {1{`RANDOM}};
  _T_257_199_1 = _RAND_797[0:0];
  _RAND_798 = {1{`RANDOM}};
  _T_257_199_2 = _RAND_798[0:0];
  _RAND_799 = {1{`RANDOM}};
  _T_257_199_3 = _RAND_799[0:0];
  _RAND_800 = {1{`RANDOM}};
  _T_257_200_0 = _RAND_800[0:0];
  _RAND_801 = {1{`RANDOM}};
  _T_257_200_1 = _RAND_801[0:0];
  _RAND_802 = {1{`RANDOM}};
  _T_257_200_2 = _RAND_802[0:0];
  _RAND_803 = {1{`RANDOM}};
  _T_257_200_3 = _RAND_803[0:0];
  _RAND_804 = {1{`RANDOM}};
  _T_257_201_0 = _RAND_804[0:0];
  _RAND_805 = {1{`RANDOM}};
  _T_257_201_1 = _RAND_805[0:0];
  _RAND_806 = {1{`RANDOM}};
  _T_257_201_2 = _RAND_806[0:0];
  _RAND_807 = {1{`RANDOM}};
  _T_257_201_3 = _RAND_807[0:0];
  _RAND_808 = {1{`RANDOM}};
  _T_257_202_0 = _RAND_808[0:0];
  _RAND_809 = {1{`RANDOM}};
  _T_257_202_1 = _RAND_809[0:0];
  _RAND_810 = {1{`RANDOM}};
  _T_257_202_2 = _RAND_810[0:0];
  _RAND_811 = {1{`RANDOM}};
  _T_257_202_3 = _RAND_811[0:0];
  _RAND_812 = {1{`RANDOM}};
  _T_257_203_0 = _RAND_812[0:0];
  _RAND_813 = {1{`RANDOM}};
  _T_257_203_1 = _RAND_813[0:0];
  _RAND_814 = {1{`RANDOM}};
  _T_257_203_2 = _RAND_814[0:0];
  _RAND_815 = {1{`RANDOM}};
  _T_257_203_3 = _RAND_815[0:0];
  _RAND_816 = {1{`RANDOM}};
  _T_257_204_0 = _RAND_816[0:0];
  _RAND_817 = {1{`RANDOM}};
  _T_257_204_1 = _RAND_817[0:0];
  _RAND_818 = {1{`RANDOM}};
  _T_257_204_2 = _RAND_818[0:0];
  _RAND_819 = {1{`RANDOM}};
  _T_257_204_3 = _RAND_819[0:0];
  _RAND_820 = {1{`RANDOM}};
  _T_257_205_0 = _RAND_820[0:0];
  _RAND_821 = {1{`RANDOM}};
  _T_257_205_1 = _RAND_821[0:0];
  _RAND_822 = {1{`RANDOM}};
  _T_257_205_2 = _RAND_822[0:0];
  _RAND_823 = {1{`RANDOM}};
  _T_257_205_3 = _RAND_823[0:0];
  _RAND_824 = {1{`RANDOM}};
  _T_257_206_0 = _RAND_824[0:0];
  _RAND_825 = {1{`RANDOM}};
  _T_257_206_1 = _RAND_825[0:0];
  _RAND_826 = {1{`RANDOM}};
  _T_257_206_2 = _RAND_826[0:0];
  _RAND_827 = {1{`RANDOM}};
  _T_257_206_3 = _RAND_827[0:0];
  _RAND_828 = {1{`RANDOM}};
  _T_257_207_0 = _RAND_828[0:0];
  _RAND_829 = {1{`RANDOM}};
  _T_257_207_1 = _RAND_829[0:0];
  _RAND_830 = {1{`RANDOM}};
  _T_257_207_2 = _RAND_830[0:0];
  _RAND_831 = {1{`RANDOM}};
  _T_257_207_3 = _RAND_831[0:0];
  _RAND_832 = {1{`RANDOM}};
  _T_257_208_0 = _RAND_832[0:0];
  _RAND_833 = {1{`RANDOM}};
  _T_257_208_1 = _RAND_833[0:0];
  _RAND_834 = {1{`RANDOM}};
  _T_257_208_2 = _RAND_834[0:0];
  _RAND_835 = {1{`RANDOM}};
  _T_257_208_3 = _RAND_835[0:0];
  _RAND_836 = {1{`RANDOM}};
  _T_257_209_0 = _RAND_836[0:0];
  _RAND_837 = {1{`RANDOM}};
  _T_257_209_1 = _RAND_837[0:0];
  _RAND_838 = {1{`RANDOM}};
  _T_257_209_2 = _RAND_838[0:0];
  _RAND_839 = {1{`RANDOM}};
  _T_257_209_3 = _RAND_839[0:0];
  _RAND_840 = {1{`RANDOM}};
  _T_257_210_0 = _RAND_840[0:0];
  _RAND_841 = {1{`RANDOM}};
  _T_257_210_1 = _RAND_841[0:0];
  _RAND_842 = {1{`RANDOM}};
  _T_257_210_2 = _RAND_842[0:0];
  _RAND_843 = {1{`RANDOM}};
  _T_257_210_3 = _RAND_843[0:0];
  _RAND_844 = {1{`RANDOM}};
  _T_257_211_0 = _RAND_844[0:0];
  _RAND_845 = {1{`RANDOM}};
  _T_257_211_1 = _RAND_845[0:0];
  _RAND_846 = {1{`RANDOM}};
  _T_257_211_2 = _RAND_846[0:0];
  _RAND_847 = {1{`RANDOM}};
  _T_257_211_3 = _RAND_847[0:0];
  _RAND_848 = {1{`RANDOM}};
  _T_257_212_0 = _RAND_848[0:0];
  _RAND_849 = {1{`RANDOM}};
  _T_257_212_1 = _RAND_849[0:0];
  _RAND_850 = {1{`RANDOM}};
  _T_257_212_2 = _RAND_850[0:0];
  _RAND_851 = {1{`RANDOM}};
  _T_257_212_3 = _RAND_851[0:0];
  _RAND_852 = {1{`RANDOM}};
  _T_257_213_0 = _RAND_852[0:0];
  _RAND_853 = {1{`RANDOM}};
  _T_257_213_1 = _RAND_853[0:0];
  _RAND_854 = {1{`RANDOM}};
  _T_257_213_2 = _RAND_854[0:0];
  _RAND_855 = {1{`RANDOM}};
  _T_257_213_3 = _RAND_855[0:0];
  _RAND_856 = {1{`RANDOM}};
  _T_257_214_0 = _RAND_856[0:0];
  _RAND_857 = {1{`RANDOM}};
  _T_257_214_1 = _RAND_857[0:0];
  _RAND_858 = {1{`RANDOM}};
  _T_257_214_2 = _RAND_858[0:0];
  _RAND_859 = {1{`RANDOM}};
  _T_257_214_3 = _RAND_859[0:0];
  _RAND_860 = {1{`RANDOM}};
  _T_257_215_0 = _RAND_860[0:0];
  _RAND_861 = {1{`RANDOM}};
  _T_257_215_1 = _RAND_861[0:0];
  _RAND_862 = {1{`RANDOM}};
  _T_257_215_2 = _RAND_862[0:0];
  _RAND_863 = {1{`RANDOM}};
  _T_257_215_3 = _RAND_863[0:0];
  _RAND_864 = {1{`RANDOM}};
  _T_257_216_0 = _RAND_864[0:0];
  _RAND_865 = {1{`RANDOM}};
  _T_257_216_1 = _RAND_865[0:0];
  _RAND_866 = {1{`RANDOM}};
  _T_257_216_2 = _RAND_866[0:0];
  _RAND_867 = {1{`RANDOM}};
  _T_257_216_3 = _RAND_867[0:0];
  _RAND_868 = {1{`RANDOM}};
  _T_257_217_0 = _RAND_868[0:0];
  _RAND_869 = {1{`RANDOM}};
  _T_257_217_1 = _RAND_869[0:0];
  _RAND_870 = {1{`RANDOM}};
  _T_257_217_2 = _RAND_870[0:0];
  _RAND_871 = {1{`RANDOM}};
  _T_257_217_3 = _RAND_871[0:0];
  _RAND_872 = {1{`RANDOM}};
  _T_257_218_0 = _RAND_872[0:0];
  _RAND_873 = {1{`RANDOM}};
  _T_257_218_1 = _RAND_873[0:0];
  _RAND_874 = {1{`RANDOM}};
  _T_257_218_2 = _RAND_874[0:0];
  _RAND_875 = {1{`RANDOM}};
  _T_257_218_3 = _RAND_875[0:0];
  _RAND_876 = {1{`RANDOM}};
  _T_257_219_0 = _RAND_876[0:0];
  _RAND_877 = {1{`RANDOM}};
  _T_257_219_1 = _RAND_877[0:0];
  _RAND_878 = {1{`RANDOM}};
  _T_257_219_2 = _RAND_878[0:0];
  _RAND_879 = {1{`RANDOM}};
  _T_257_219_3 = _RAND_879[0:0];
  _RAND_880 = {1{`RANDOM}};
  _T_257_220_0 = _RAND_880[0:0];
  _RAND_881 = {1{`RANDOM}};
  _T_257_220_1 = _RAND_881[0:0];
  _RAND_882 = {1{`RANDOM}};
  _T_257_220_2 = _RAND_882[0:0];
  _RAND_883 = {1{`RANDOM}};
  _T_257_220_3 = _RAND_883[0:0];
  _RAND_884 = {1{`RANDOM}};
  _T_257_221_0 = _RAND_884[0:0];
  _RAND_885 = {1{`RANDOM}};
  _T_257_221_1 = _RAND_885[0:0];
  _RAND_886 = {1{`RANDOM}};
  _T_257_221_2 = _RAND_886[0:0];
  _RAND_887 = {1{`RANDOM}};
  _T_257_221_3 = _RAND_887[0:0];
  _RAND_888 = {1{`RANDOM}};
  _T_257_222_0 = _RAND_888[0:0];
  _RAND_889 = {1{`RANDOM}};
  _T_257_222_1 = _RAND_889[0:0];
  _RAND_890 = {1{`RANDOM}};
  _T_257_222_2 = _RAND_890[0:0];
  _RAND_891 = {1{`RANDOM}};
  _T_257_222_3 = _RAND_891[0:0];
  _RAND_892 = {1{`RANDOM}};
  _T_257_223_0 = _RAND_892[0:0];
  _RAND_893 = {1{`RANDOM}};
  _T_257_223_1 = _RAND_893[0:0];
  _RAND_894 = {1{`RANDOM}};
  _T_257_223_2 = _RAND_894[0:0];
  _RAND_895 = {1{`RANDOM}};
  _T_257_223_3 = _RAND_895[0:0];
  _RAND_896 = {1{`RANDOM}};
  _T_257_224_0 = _RAND_896[0:0];
  _RAND_897 = {1{`RANDOM}};
  _T_257_224_1 = _RAND_897[0:0];
  _RAND_898 = {1{`RANDOM}};
  _T_257_224_2 = _RAND_898[0:0];
  _RAND_899 = {1{`RANDOM}};
  _T_257_224_3 = _RAND_899[0:0];
  _RAND_900 = {1{`RANDOM}};
  _T_257_225_0 = _RAND_900[0:0];
  _RAND_901 = {1{`RANDOM}};
  _T_257_225_1 = _RAND_901[0:0];
  _RAND_902 = {1{`RANDOM}};
  _T_257_225_2 = _RAND_902[0:0];
  _RAND_903 = {1{`RANDOM}};
  _T_257_225_3 = _RAND_903[0:0];
  _RAND_904 = {1{`RANDOM}};
  _T_257_226_0 = _RAND_904[0:0];
  _RAND_905 = {1{`RANDOM}};
  _T_257_226_1 = _RAND_905[0:0];
  _RAND_906 = {1{`RANDOM}};
  _T_257_226_2 = _RAND_906[0:0];
  _RAND_907 = {1{`RANDOM}};
  _T_257_226_3 = _RAND_907[0:0];
  _RAND_908 = {1{`RANDOM}};
  _T_257_227_0 = _RAND_908[0:0];
  _RAND_909 = {1{`RANDOM}};
  _T_257_227_1 = _RAND_909[0:0];
  _RAND_910 = {1{`RANDOM}};
  _T_257_227_2 = _RAND_910[0:0];
  _RAND_911 = {1{`RANDOM}};
  _T_257_227_3 = _RAND_911[0:0];
  _RAND_912 = {1{`RANDOM}};
  _T_257_228_0 = _RAND_912[0:0];
  _RAND_913 = {1{`RANDOM}};
  _T_257_228_1 = _RAND_913[0:0];
  _RAND_914 = {1{`RANDOM}};
  _T_257_228_2 = _RAND_914[0:0];
  _RAND_915 = {1{`RANDOM}};
  _T_257_228_3 = _RAND_915[0:0];
  _RAND_916 = {1{`RANDOM}};
  _T_257_229_0 = _RAND_916[0:0];
  _RAND_917 = {1{`RANDOM}};
  _T_257_229_1 = _RAND_917[0:0];
  _RAND_918 = {1{`RANDOM}};
  _T_257_229_2 = _RAND_918[0:0];
  _RAND_919 = {1{`RANDOM}};
  _T_257_229_3 = _RAND_919[0:0];
  _RAND_920 = {1{`RANDOM}};
  _T_257_230_0 = _RAND_920[0:0];
  _RAND_921 = {1{`RANDOM}};
  _T_257_230_1 = _RAND_921[0:0];
  _RAND_922 = {1{`RANDOM}};
  _T_257_230_2 = _RAND_922[0:0];
  _RAND_923 = {1{`RANDOM}};
  _T_257_230_3 = _RAND_923[0:0];
  _RAND_924 = {1{`RANDOM}};
  _T_257_231_0 = _RAND_924[0:0];
  _RAND_925 = {1{`RANDOM}};
  _T_257_231_1 = _RAND_925[0:0];
  _RAND_926 = {1{`RANDOM}};
  _T_257_231_2 = _RAND_926[0:0];
  _RAND_927 = {1{`RANDOM}};
  _T_257_231_3 = _RAND_927[0:0];
  _RAND_928 = {1{`RANDOM}};
  _T_257_232_0 = _RAND_928[0:0];
  _RAND_929 = {1{`RANDOM}};
  _T_257_232_1 = _RAND_929[0:0];
  _RAND_930 = {1{`RANDOM}};
  _T_257_232_2 = _RAND_930[0:0];
  _RAND_931 = {1{`RANDOM}};
  _T_257_232_3 = _RAND_931[0:0];
  _RAND_932 = {1{`RANDOM}};
  _T_257_233_0 = _RAND_932[0:0];
  _RAND_933 = {1{`RANDOM}};
  _T_257_233_1 = _RAND_933[0:0];
  _RAND_934 = {1{`RANDOM}};
  _T_257_233_2 = _RAND_934[0:0];
  _RAND_935 = {1{`RANDOM}};
  _T_257_233_3 = _RAND_935[0:0];
  _RAND_936 = {1{`RANDOM}};
  _T_257_234_0 = _RAND_936[0:0];
  _RAND_937 = {1{`RANDOM}};
  _T_257_234_1 = _RAND_937[0:0];
  _RAND_938 = {1{`RANDOM}};
  _T_257_234_2 = _RAND_938[0:0];
  _RAND_939 = {1{`RANDOM}};
  _T_257_234_3 = _RAND_939[0:0];
  _RAND_940 = {1{`RANDOM}};
  _T_257_235_0 = _RAND_940[0:0];
  _RAND_941 = {1{`RANDOM}};
  _T_257_235_1 = _RAND_941[0:0];
  _RAND_942 = {1{`RANDOM}};
  _T_257_235_2 = _RAND_942[0:0];
  _RAND_943 = {1{`RANDOM}};
  _T_257_235_3 = _RAND_943[0:0];
  _RAND_944 = {1{`RANDOM}};
  _T_257_236_0 = _RAND_944[0:0];
  _RAND_945 = {1{`RANDOM}};
  _T_257_236_1 = _RAND_945[0:0];
  _RAND_946 = {1{`RANDOM}};
  _T_257_236_2 = _RAND_946[0:0];
  _RAND_947 = {1{`RANDOM}};
  _T_257_236_3 = _RAND_947[0:0];
  _RAND_948 = {1{`RANDOM}};
  _T_257_237_0 = _RAND_948[0:0];
  _RAND_949 = {1{`RANDOM}};
  _T_257_237_1 = _RAND_949[0:0];
  _RAND_950 = {1{`RANDOM}};
  _T_257_237_2 = _RAND_950[0:0];
  _RAND_951 = {1{`RANDOM}};
  _T_257_237_3 = _RAND_951[0:0];
  _RAND_952 = {1{`RANDOM}};
  _T_257_238_0 = _RAND_952[0:0];
  _RAND_953 = {1{`RANDOM}};
  _T_257_238_1 = _RAND_953[0:0];
  _RAND_954 = {1{`RANDOM}};
  _T_257_238_2 = _RAND_954[0:0];
  _RAND_955 = {1{`RANDOM}};
  _T_257_238_3 = _RAND_955[0:0];
  _RAND_956 = {1{`RANDOM}};
  _T_257_239_0 = _RAND_956[0:0];
  _RAND_957 = {1{`RANDOM}};
  _T_257_239_1 = _RAND_957[0:0];
  _RAND_958 = {1{`RANDOM}};
  _T_257_239_2 = _RAND_958[0:0];
  _RAND_959 = {1{`RANDOM}};
  _T_257_239_3 = _RAND_959[0:0];
  _RAND_960 = {1{`RANDOM}};
  _T_257_240_0 = _RAND_960[0:0];
  _RAND_961 = {1{`RANDOM}};
  _T_257_240_1 = _RAND_961[0:0];
  _RAND_962 = {1{`RANDOM}};
  _T_257_240_2 = _RAND_962[0:0];
  _RAND_963 = {1{`RANDOM}};
  _T_257_240_3 = _RAND_963[0:0];
  _RAND_964 = {1{`RANDOM}};
  _T_257_241_0 = _RAND_964[0:0];
  _RAND_965 = {1{`RANDOM}};
  _T_257_241_1 = _RAND_965[0:0];
  _RAND_966 = {1{`RANDOM}};
  _T_257_241_2 = _RAND_966[0:0];
  _RAND_967 = {1{`RANDOM}};
  _T_257_241_3 = _RAND_967[0:0];
  _RAND_968 = {1{`RANDOM}};
  _T_257_242_0 = _RAND_968[0:0];
  _RAND_969 = {1{`RANDOM}};
  _T_257_242_1 = _RAND_969[0:0];
  _RAND_970 = {1{`RANDOM}};
  _T_257_242_2 = _RAND_970[0:0];
  _RAND_971 = {1{`RANDOM}};
  _T_257_242_3 = _RAND_971[0:0];
  _RAND_972 = {1{`RANDOM}};
  _T_257_243_0 = _RAND_972[0:0];
  _RAND_973 = {1{`RANDOM}};
  _T_257_243_1 = _RAND_973[0:0];
  _RAND_974 = {1{`RANDOM}};
  _T_257_243_2 = _RAND_974[0:0];
  _RAND_975 = {1{`RANDOM}};
  _T_257_243_3 = _RAND_975[0:0];
  _RAND_976 = {1{`RANDOM}};
  _T_257_244_0 = _RAND_976[0:0];
  _RAND_977 = {1{`RANDOM}};
  _T_257_244_1 = _RAND_977[0:0];
  _RAND_978 = {1{`RANDOM}};
  _T_257_244_2 = _RAND_978[0:0];
  _RAND_979 = {1{`RANDOM}};
  _T_257_244_3 = _RAND_979[0:0];
  _RAND_980 = {1{`RANDOM}};
  _T_257_245_0 = _RAND_980[0:0];
  _RAND_981 = {1{`RANDOM}};
  _T_257_245_1 = _RAND_981[0:0];
  _RAND_982 = {1{`RANDOM}};
  _T_257_245_2 = _RAND_982[0:0];
  _RAND_983 = {1{`RANDOM}};
  _T_257_245_3 = _RAND_983[0:0];
  _RAND_984 = {1{`RANDOM}};
  _T_257_246_0 = _RAND_984[0:0];
  _RAND_985 = {1{`RANDOM}};
  _T_257_246_1 = _RAND_985[0:0];
  _RAND_986 = {1{`RANDOM}};
  _T_257_246_2 = _RAND_986[0:0];
  _RAND_987 = {1{`RANDOM}};
  _T_257_246_3 = _RAND_987[0:0];
  _RAND_988 = {1{`RANDOM}};
  _T_257_247_0 = _RAND_988[0:0];
  _RAND_989 = {1{`RANDOM}};
  _T_257_247_1 = _RAND_989[0:0];
  _RAND_990 = {1{`RANDOM}};
  _T_257_247_2 = _RAND_990[0:0];
  _RAND_991 = {1{`RANDOM}};
  _T_257_247_3 = _RAND_991[0:0];
  _RAND_992 = {1{`RANDOM}};
  _T_257_248_0 = _RAND_992[0:0];
  _RAND_993 = {1{`RANDOM}};
  _T_257_248_1 = _RAND_993[0:0];
  _RAND_994 = {1{`RANDOM}};
  _T_257_248_2 = _RAND_994[0:0];
  _RAND_995 = {1{`RANDOM}};
  _T_257_248_3 = _RAND_995[0:0];
  _RAND_996 = {1{`RANDOM}};
  _T_257_249_0 = _RAND_996[0:0];
  _RAND_997 = {1{`RANDOM}};
  _T_257_249_1 = _RAND_997[0:0];
  _RAND_998 = {1{`RANDOM}};
  _T_257_249_2 = _RAND_998[0:0];
  _RAND_999 = {1{`RANDOM}};
  _T_257_249_3 = _RAND_999[0:0];
  _RAND_1000 = {1{`RANDOM}};
  _T_257_250_0 = _RAND_1000[0:0];
  _RAND_1001 = {1{`RANDOM}};
  _T_257_250_1 = _RAND_1001[0:0];
  _RAND_1002 = {1{`RANDOM}};
  _T_257_250_2 = _RAND_1002[0:0];
  _RAND_1003 = {1{`RANDOM}};
  _T_257_250_3 = _RAND_1003[0:0];
  _RAND_1004 = {1{`RANDOM}};
  _T_257_251_0 = _RAND_1004[0:0];
  _RAND_1005 = {1{`RANDOM}};
  _T_257_251_1 = _RAND_1005[0:0];
  _RAND_1006 = {1{`RANDOM}};
  _T_257_251_2 = _RAND_1006[0:0];
  _RAND_1007 = {1{`RANDOM}};
  _T_257_251_3 = _RAND_1007[0:0];
  _RAND_1008 = {1{`RANDOM}};
  _T_257_252_0 = _RAND_1008[0:0];
  _RAND_1009 = {1{`RANDOM}};
  _T_257_252_1 = _RAND_1009[0:0];
  _RAND_1010 = {1{`RANDOM}};
  _T_257_252_2 = _RAND_1010[0:0];
  _RAND_1011 = {1{`RANDOM}};
  _T_257_252_3 = _RAND_1011[0:0];
  _RAND_1012 = {1{`RANDOM}};
  _T_257_253_0 = _RAND_1012[0:0];
  _RAND_1013 = {1{`RANDOM}};
  _T_257_253_1 = _RAND_1013[0:0];
  _RAND_1014 = {1{`RANDOM}};
  _T_257_253_2 = _RAND_1014[0:0];
  _RAND_1015 = {1{`RANDOM}};
  _T_257_253_3 = _RAND_1015[0:0];
  _RAND_1016 = {1{`RANDOM}};
  _T_257_254_0 = _RAND_1016[0:0];
  _RAND_1017 = {1{`RANDOM}};
  _T_257_254_1 = _RAND_1017[0:0];
  _RAND_1018 = {1{`RANDOM}};
  _T_257_254_2 = _RAND_1018[0:0];
  _RAND_1019 = {1{`RANDOM}};
  _T_257_254_3 = _RAND_1019[0:0];
  _RAND_1020 = {1{`RANDOM}};
  _T_257_255_0 = _RAND_1020[0:0];
  _RAND_1021 = {1{`RANDOM}};
  _T_257_255_1 = _RAND_1021[0:0];
  _RAND_1022 = {1{`RANDOM}};
  _T_257_255_2 = _RAND_1022[0:0];
  _RAND_1023 = {1{`RANDOM}};
  _T_257_255_3 = _RAND_1023[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      _T_257_0_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h0 == io_fetchQuery_index) begin
        if (_T_300) begin
          _T_257_0_0 <= _GEN_4108;
        end else begin
          _T_257_0_0 <= _GEN_2052;
        end
      end
    end
    if (reset) begin
      _T_257_0_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h0 == io_fetchQuery_index) begin
        if (_T_300) begin
          _T_257_0_1 <= _GEN_4109;
        end else begin
          _T_257_0_1 <= _GEN_2053;
        end
      end
    end
    if (reset) begin
      _T_257_0_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h0 == io_fetchQuery_index) begin
        if (_T_300) begin
          _T_257_0_2 <= _GEN_4110;
        end else begin
          _T_257_0_2 <= _GEN_2054;
        end
      end
    end
    if (reset) begin
      _T_257_0_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h0 == io_fetchQuery_index) begin
        if (_T_300) begin
          _T_257_0_3 <= _GEN_4111;
        end else begin
          _T_257_0_3 <= _GEN_2055;
        end
      end
    end
    if (reset) begin
      _T_257_1_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h1 == io_fetchQuery_index) begin
        if (_T_300) begin
          _T_257_1_0 <= _GEN_4108;
        end else begin
          _T_257_1_0 <= _GEN_2052;
        end
      end
    end
    if (reset) begin
      _T_257_1_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h1 == io_fetchQuery_index) begin
        if (_T_300) begin
          _T_257_1_1 <= _GEN_4109;
        end else begin
          _T_257_1_1 <= _GEN_2053;
        end
      end
    end
    if (reset) begin
      _T_257_1_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h1 == io_fetchQuery_index) begin
        if (_T_300) begin
          _T_257_1_2 <= _GEN_4110;
        end else begin
          _T_257_1_2 <= _GEN_2054;
        end
      end
    end
    if (reset) begin
      _T_257_1_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h1 == io_fetchQuery_index) begin
        if (_T_300) begin
          _T_257_1_3 <= _GEN_4111;
        end else begin
          _T_257_1_3 <= _GEN_2055;
        end
      end
    end
    if (reset) begin
      _T_257_2_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h2 == io_fetchQuery_index) begin
        if (_T_300) begin
          _T_257_2_0 <= _GEN_4108;
        end else begin
          _T_257_2_0 <= _GEN_2052;
        end
      end
    end
    if (reset) begin
      _T_257_2_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h2 == io_fetchQuery_index) begin
        if (_T_300) begin
          _T_257_2_1 <= _GEN_4109;
        end else begin
          _T_257_2_1 <= _GEN_2053;
        end
      end
    end
    if (reset) begin
      _T_257_2_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h2 == io_fetchQuery_index) begin
        if (_T_300) begin
          _T_257_2_2 <= _GEN_4110;
        end else begin
          _T_257_2_2 <= _GEN_2054;
        end
      end
    end
    if (reset) begin
      _T_257_2_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h2 == io_fetchQuery_index) begin
        if (_T_300) begin
          _T_257_2_3 <= _GEN_4111;
        end else begin
          _T_257_2_3 <= _GEN_2055;
        end
      end
    end
    if (reset) begin
      _T_257_3_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h3 == io_fetchQuery_index) begin
        if (_T_300) begin
          _T_257_3_0 <= _GEN_4108;
        end else begin
          _T_257_3_0 <= _GEN_2052;
        end
      end
    end
    if (reset) begin
      _T_257_3_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h3 == io_fetchQuery_index) begin
        if (_T_300) begin
          _T_257_3_1 <= _GEN_4109;
        end else begin
          _T_257_3_1 <= _GEN_2053;
        end
      end
    end
    if (reset) begin
      _T_257_3_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h3 == io_fetchQuery_index) begin
        if (_T_300) begin
          _T_257_3_2 <= _GEN_4110;
        end else begin
          _T_257_3_2 <= _GEN_2054;
        end
      end
    end
    if (reset) begin
      _T_257_3_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h3 == io_fetchQuery_index) begin
        if (_T_300) begin
          _T_257_3_3 <= _GEN_4111;
        end else begin
          _T_257_3_3 <= _GEN_2055;
        end
      end
    end
    if (reset) begin
      _T_257_4_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h4 == io_fetchQuery_index) begin
        _T_257_4_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_4_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h4 == io_fetchQuery_index) begin
        _T_257_4_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_4_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h4 == io_fetchQuery_index) begin
        _T_257_4_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_4_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h4 == io_fetchQuery_index) begin
        _T_257_4_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_5_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h5 == io_fetchQuery_index) begin
        _T_257_5_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_5_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h5 == io_fetchQuery_index) begin
        _T_257_5_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_5_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h5 == io_fetchQuery_index) begin
        _T_257_5_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_5_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h5 == io_fetchQuery_index) begin
        _T_257_5_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_6_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h6 == io_fetchQuery_index) begin
        _T_257_6_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_6_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h6 == io_fetchQuery_index) begin
        _T_257_6_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_6_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h6 == io_fetchQuery_index) begin
        _T_257_6_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_6_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h6 == io_fetchQuery_index) begin
        _T_257_6_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_7_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h7 == io_fetchQuery_index) begin
        _T_257_7_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_7_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h7 == io_fetchQuery_index) begin
        _T_257_7_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_7_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h7 == io_fetchQuery_index) begin
        _T_257_7_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_7_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h7 == io_fetchQuery_index) begin
        _T_257_7_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_8_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h8 == io_fetchQuery_index) begin
        _T_257_8_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_8_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h8 == io_fetchQuery_index) begin
        _T_257_8_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_8_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h8 == io_fetchQuery_index) begin
        _T_257_8_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_8_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h8 == io_fetchQuery_index) begin
        _T_257_8_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_9_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h9 == io_fetchQuery_index) begin
        _T_257_9_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_9_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h9 == io_fetchQuery_index) begin
        _T_257_9_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_9_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h9 == io_fetchQuery_index) begin
        _T_257_9_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_9_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h9 == io_fetchQuery_index) begin
        _T_257_9_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_10_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'ha == io_fetchQuery_index) begin
        _T_257_10_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_10_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'ha == io_fetchQuery_index) begin
        _T_257_10_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_10_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'ha == io_fetchQuery_index) begin
        _T_257_10_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_10_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'ha == io_fetchQuery_index) begin
        _T_257_10_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_11_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hb == io_fetchQuery_index) begin
        _T_257_11_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_11_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hb == io_fetchQuery_index) begin
        _T_257_11_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_11_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hb == io_fetchQuery_index) begin
        _T_257_11_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_11_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hb == io_fetchQuery_index) begin
        _T_257_11_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_12_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hc == io_fetchQuery_index) begin
        _T_257_12_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_12_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hc == io_fetchQuery_index) begin
        _T_257_12_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_12_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hc == io_fetchQuery_index) begin
        _T_257_12_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_12_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hc == io_fetchQuery_index) begin
        _T_257_12_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_13_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hd == io_fetchQuery_index) begin
        _T_257_13_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_13_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hd == io_fetchQuery_index) begin
        _T_257_13_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_13_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hd == io_fetchQuery_index) begin
        _T_257_13_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_13_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hd == io_fetchQuery_index) begin
        _T_257_13_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_14_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'he == io_fetchQuery_index) begin
        _T_257_14_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_14_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'he == io_fetchQuery_index) begin
        _T_257_14_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_14_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'he == io_fetchQuery_index) begin
        _T_257_14_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_14_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'he == io_fetchQuery_index) begin
        _T_257_14_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_15_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hf == io_fetchQuery_index) begin
        _T_257_15_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_15_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hf == io_fetchQuery_index) begin
        _T_257_15_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_15_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hf == io_fetchQuery_index) begin
        _T_257_15_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_15_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hf == io_fetchQuery_index) begin
        _T_257_15_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_16_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h10 == io_fetchQuery_index) begin
        _T_257_16_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_16_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h10 == io_fetchQuery_index) begin
        _T_257_16_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_16_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h10 == io_fetchQuery_index) begin
        _T_257_16_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_16_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h10 == io_fetchQuery_index) begin
        _T_257_16_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_17_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h11 == io_fetchQuery_index) begin
        _T_257_17_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_17_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h11 == io_fetchQuery_index) begin
        _T_257_17_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_17_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h11 == io_fetchQuery_index) begin
        _T_257_17_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_17_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h11 == io_fetchQuery_index) begin
        _T_257_17_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_18_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h12 == io_fetchQuery_index) begin
        _T_257_18_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_18_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h12 == io_fetchQuery_index) begin
        _T_257_18_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_18_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h12 == io_fetchQuery_index) begin
        _T_257_18_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_18_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h12 == io_fetchQuery_index) begin
        _T_257_18_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_19_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h13 == io_fetchQuery_index) begin
        _T_257_19_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_19_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h13 == io_fetchQuery_index) begin
        _T_257_19_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_19_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h13 == io_fetchQuery_index) begin
        _T_257_19_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_19_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h13 == io_fetchQuery_index) begin
        _T_257_19_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_20_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h14 == io_fetchQuery_index) begin
        _T_257_20_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_20_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h14 == io_fetchQuery_index) begin
        _T_257_20_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_20_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h14 == io_fetchQuery_index) begin
        _T_257_20_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_20_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h14 == io_fetchQuery_index) begin
        _T_257_20_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_21_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h15 == io_fetchQuery_index) begin
        _T_257_21_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_21_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h15 == io_fetchQuery_index) begin
        _T_257_21_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_21_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h15 == io_fetchQuery_index) begin
        _T_257_21_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_21_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h15 == io_fetchQuery_index) begin
        _T_257_21_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_22_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h16 == io_fetchQuery_index) begin
        _T_257_22_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_22_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h16 == io_fetchQuery_index) begin
        _T_257_22_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_22_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h16 == io_fetchQuery_index) begin
        _T_257_22_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_22_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h16 == io_fetchQuery_index) begin
        _T_257_22_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_23_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h17 == io_fetchQuery_index) begin
        _T_257_23_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_23_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h17 == io_fetchQuery_index) begin
        _T_257_23_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_23_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h17 == io_fetchQuery_index) begin
        _T_257_23_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_23_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h17 == io_fetchQuery_index) begin
        _T_257_23_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_24_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h18 == io_fetchQuery_index) begin
        _T_257_24_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_24_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h18 == io_fetchQuery_index) begin
        _T_257_24_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_24_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h18 == io_fetchQuery_index) begin
        _T_257_24_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_24_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h18 == io_fetchQuery_index) begin
        _T_257_24_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_25_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h19 == io_fetchQuery_index) begin
        _T_257_25_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_25_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h19 == io_fetchQuery_index) begin
        _T_257_25_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_25_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h19 == io_fetchQuery_index) begin
        _T_257_25_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_25_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h19 == io_fetchQuery_index) begin
        _T_257_25_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_26_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h1a == io_fetchQuery_index) begin
        _T_257_26_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_26_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h1a == io_fetchQuery_index) begin
        _T_257_26_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_26_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h1a == io_fetchQuery_index) begin
        _T_257_26_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_26_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h1a == io_fetchQuery_index) begin
        _T_257_26_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_27_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h1b == io_fetchQuery_index) begin
        _T_257_27_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_27_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h1b == io_fetchQuery_index) begin
        _T_257_27_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_27_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h1b == io_fetchQuery_index) begin
        _T_257_27_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_27_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h1b == io_fetchQuery_index) begin
        _T_257_27_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_28_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h1c == io_fetchQuery_index) begin
        _T_257_28_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_28_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h1c == io_fetchQuery_index) begin
        _T_257_28_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_28_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h1c == io_fetchQuery_index) begin
        _T_257_28_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_28_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h1c == io_fetchQuery_index) begin
        _T_257_28_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_29_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h1d == io_fetchQuery_index) begin
        _T_257_29_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_29_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h1d == io_fetchQuery_index) begin
        _T_257_29_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_29_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h1d == io_fetchQuery_index) begin
        _T_257_29_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_29_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h1d == io_fetchQuery_index) begin
        _T_257_29_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_30_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h1e == io_fetchQuery_index) begin
        _T_257_30_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_30_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h1e == io_fetchQuery_index) begin
        _T_257_30_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_30_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h1e == io_fetchQuery_index) begin
        _T_257_30_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_30_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h1e == io_fetchQuery_index) begin
        _T_257_30_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_31_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h1f == io_fetchQuery_index) begin
        _T_257_31_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_31_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h1f == io_fetchQuery_index) begin
        _T_257_31_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_31_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h1f == io_fetchQuery_index) begin
        _T_257_31_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_31_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h1f == io_fetchQuery_index) begin
        _T_257_31_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_32_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h20 == io_fetchQuery_index) begin
        _T_257_32_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_32_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h20 == io_fetchQuery_index) begin
        _T_257_32_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_32_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h20 == io_fetchQuery_index) begin
        _T_257_32_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_32_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h20 == io_fetchQuery_index) begin
        _T_257_32_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_33_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h21 == io_fetchQuery_index) begin
        _T_257_33_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_33_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h21 == io_fetchQuery_index) begin
        _T_257_33_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_33_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h21 == io_fetchQuery_index) begin
        _T_257_33_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_33_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h21 == io_fetchQuery_index) begin
        _T_257_33_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_34_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h22 == io_fetchQuery_index) begin
        _T_257_34_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_34_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h22 == io_fetchQuery_index) begin
        _T_257_34_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_34_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h22 == io_fetchQuery_index) begin
        _T_257_34_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_34_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h22 == io_fetchQuery_index) begin
        _T_257_34_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_35_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h23 == io_fetchQuery_index) begin
        _T_257_35_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_35_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h23 == io_fetchQuery_index) begin
        _T_257_35_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_35_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h23 == io_fetchQuery_index) begin
        _T_257_35_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_35_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h23 == io_fetchQuery_index) begin
        _T_257_35_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_36_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h24 == io_fetchQuery_index) begin
        _T_257_36_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_36_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h24 == io_fetchQuery_index) begin
        _T_257_36_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_36_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h24 == io_fetchQuery_index) begin
        _T_257_36_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_36_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h24 == io_fetchQuery_index) begin
        _T_257_36_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_37_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h25 == io_fetchQuery_index) begin
        _T_257_37_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_37_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h25 == io_fetchQuery_index) begin
        _T_257_37_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_37_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h25 == io_fetchQuery_index) begin
        _T_257_37_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_37_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h25 == io_fetchQuery_index) begin
        _T_257_37_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_38_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h26 == io_fetchQuery_index) begin
        _T_257_38_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_38_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h26 == io_fetchQuery_index) begin
        _T_257_38_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_38_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h26 == io_fetchQuery_index) begin
        _T_257_38_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_38_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h26 == io_fetchQuery_index) begin
        _T_257_38_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_39_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h27 == io_fetchQuery_index) begin
        _T_257_39_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_39_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h27 == io_fetchQuery_index) begin
        _T_257_39_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_39_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h27 == io_fetchQuery_index) begin
        _T_257_39_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_39_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h27 == io_fetchQuery_index) begin
        _T_257_39_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_40_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h28 == io_fetchQuery_index) begin
        _T_257_40_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_40_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h28 == io_fetchQuery_index) begin
        _T_257_40_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_40_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h28 == io_fetchQuery_index) begin
        _T_257_40_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_40_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h28 == io_fetchQuery_index) begin
        _T_257_40_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_41_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h29 == io_fetchQuery_index) begin
        _T_257_41_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_41_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h29 == io_fetchQuery_index) begin
        _T_257_41_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_41_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h29 == io_fetchQuery_index) begin
        _T_257_41_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_41_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h29 == io_fetchQuery_index) begin
        _T_257_41_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_42_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h2a == io_fetchQuery_index) begin
        _T_257_42_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_42_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h2a == io_fetchQuery_index) begin
        _T_257_42_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_42_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h2a == io_fetchQuery_index) begin
        _T_257_42_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_42_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h2a == io_fetchQuery_index) begin
        _T_257_42_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_43_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h2b == io_fetchQuery_index) begin
        _T_257_43_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_43_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h2b == io_fetchQuery_index) begin
        _T_257_43_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_43_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h2b == io_fetchQuery_index) begin
        _T_257_43_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_43_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h2b == io_fetchQuery_index) begin
        _T_257_43_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_44_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h2c == io_fetchQuery_index) begin
        _T_257_44_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_44_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h2c == io_fetchQuery_index) begin
        _T_257_44_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_44_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h2c == io_fetchQuery_index) begin
        _T_257_44_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_44_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h2c == io_fetchQuery_index) begin
        _T_257_44_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_45_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h2d == io_fetchQuery_index) begin
        _T_257_45_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_45_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h2d == io_fetchQuery_index) begin
        _T_257_45_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_45_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h2d == io_fetchQuery_index) begin
        _T_257_45_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_45_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h2d == io_fetchQuery_index) begin
        _T_257_45_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_46_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h2e == io_fetchQuery_index) begin
        _T_257_46_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_46_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h2e == io_fetchQuery_index) begin
        _T_257_46_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_46_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h2e == io_fetchQuery_index) begin
        _T_257_46_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_46_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h2e == io_fetchQuery_index) begin
        _T_257_46_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_47_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h2f == io_fetchQuery_index) begin
        _T_257_47_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_47_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h2f == io_fetchQuery_index) begin
        _T_257_47_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_47_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h2f == io_fetchQuery_index) begin
        _T_257_47_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_47_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h2f == io_fetchQuery_index) begin
        _T_257_47_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_48_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h30 == io_fetchQuery_index) begin
        _T_257_48_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_48_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h30 == io_fetchQuery_index) begin
        _T_257_48_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_48_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h30 == io_fetchQuery_index) begin
        _T_257_48_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_48_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h30 == io_fetchQuery_index) begin
        _T_257_48_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_49_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h31 == io_fetchQuery_index) begin
        _T_257_49_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_49_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h31 == io_fetchQuery_index) begin
        _T_257_49_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_49_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h31 == io_fetchQuery_index) begin
        _T_257_49_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_49_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h31 == io_fetchQuery_index) begin
        _T_257_49_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_50_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h32 == io_fetchQuery_index) begin
        _T_257_50_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_50_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h32 == io_fetchQuery_index) begin
        _T_257_50_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_50_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h32 == io_fetchQuery_index) begin
        _T_257_50_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_50_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h32 == io_fetchQuery_index) begin
        _T_257_50_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_51_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h33 == io_fetchQuery_index) begin
        _T_257_51_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_51_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h33 == io_fetchQuery_index) begin
        _T_257_51_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_51_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h33 == io_fetchQuery_index) begin
        _T_257_51_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_51_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h33 == io_fetchQuery_index) begin
        _T_257_51_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_52_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h34 == io_fetchQuery_index) begin
        _T_257_52_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_52_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h34 == io_fetchQuery_index) begin
        _T_257_52_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_52_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h34 == io_fetchQuery_index) begin
        _T_257_52_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_52_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h34 == io_fetchQuery_index) begin
        _T_257_52_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_53_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h35 == io_fetchQuery_index) begin
        _T_257_53_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_53_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h35 == io_fetchQuery_index) begin
        _T_257_53_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_53_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h35 == io_fetchQuery_index) begin
        _T_257_53_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_53_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h35 == io_fetchQuery_index) begin
        _T_257_53_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_54_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h36 == io_fetchQuery_index) begin
        _T_257_54_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_54_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h36 == io_fetchQuery_index) begin
        _T_257_54_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_54_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h36 == io_fetchQuery_index) begin
        _T_257_54_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_54_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h36 == io_fetchQuery_index) begin
        _T_257_54_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_55_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h37 == io_fetchQuery_index) begin
        _T_257_55_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_55_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h37 == io_fetchQuery_index) begin
        _T_257_55_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_55_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h37 == io_fetchQuery_index) begin
        _T_257_55_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_55_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h37 == io_fetchQuery_index) begin
        _T_257_55_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_56_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h38 == io_fetchQuery_index) begin
        _T_257_56_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_56_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h38 == io_fetchQuery_index) begin
        _T_257_56_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_56_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h38 == io_fetchQuery_index) begin
        _T_257_56_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_56_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h38 == io_fetchQuery_index) begin
        _T_257_56_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_57_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h39 == io_fetchQuery_index) begin
        _T_257_57_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_57_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h39 == io_fetchQuery_index) begin
        _T_257_57_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_57_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h39 == io_fetchQuery_index) begin
        _T_257_57_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_57_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h39 == io_fetchQuery_index) begin
        _T_257_57_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_58_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h3a == io_fetchQuery_index) begin
        _T_257_58_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_58_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h3a == io_fetchQuery_index) begin
        _T_257_58_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_58_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h3a == io_fetchQuery_index) begin
        _T_257_58_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_58_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h3a == io_fetchQuery_index) begin
        _T_257_58_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_59_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h3b == io_fetchQuery_index) begin
        _T_257_59_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_59_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h3b == io_fetchQuery_index) begin
        _T_257_59_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_59_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h3b == io_fetchQuery_index) begin
        _T_257_59_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_59_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h3b == io_fetchQuery_index) begin
        _T_257_59_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_60_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h3c == io_fetchQuery_index) begin
        _T_257_60_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_60_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h3c == io_fetchQuery_index) begin
        _T_257_60_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_60_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h3c == io_fetchQuery_index) begin
        _T_257_60_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_60_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h3c == io_fetchQuery_index) begin
        _T_257_60_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_61_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h3d == io_fetchQuery_index) begin
        _T_257_61_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_61_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h3d == io_fetchQuery_index) begin
        _T_257_61_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_61_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h3d == io_fetchQuery_index) begin
        _T_257_61_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_61_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h3d == io_fetchQuery_index) begin
        _T_257_61_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_62_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h3e == io_fetchQuery_index) begin
        _T_257_62_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_62_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h3e == io_fetchQuery_index) begin
        _T_257_62_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_62_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h3e == io_fetchQuery_index) begin
        _T_257_62_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_62_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h3e == io_fetchQuery_index) begin
        _T_257_62_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_63_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h3f == io_fetchQuery_index) begin
        _T_257_63_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_63_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h3f == io_fetchQuery_index) begin
        _T_257_63_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_63_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h3f == io_fetchQuery_index) begin
        _T_257_63_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_63_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h3f == io_fetchQuery_index) begin
        _T_257_63_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_64_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h40 == io_fetchQuery_index) begin
        _T_257_64_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_64_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h40 == io_fetchQuery_index) begin
        _T_257_64_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_64_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h40 == io_fetchQuery_index) begin
        _T_257_64_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_64_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h40 == io_fetchQuery_index) begin
        _T_257_64_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_65_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h41 == io_fetchQuery_index) begin
        _T_257_65_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_65_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h41 == io_fetchQuery_index) begin
        _T_257_65_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_65_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h41 == io_fetchQuery_index) begin
        _T_257_65_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_65_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h41 == io_fetchQuery_index) begin
        _T_257_65_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_66_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h42 == io_fetchQuery_index) begin
        _T_257_66_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_66_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h42 == io_fetchQuery_index) begin
        _T_257_66_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_66_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h42 == io_fetchQuery_index) begin
        _T_257_66_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_66_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h42 == io_fetchQuery_index) begin
        _T_257_66_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_67_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h43 == io_fetchQuery_index) begin
        _T_257_67_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_67_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h43 == io_fetchQuery_index) begin
        _T_257_67_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_67_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h43 == io_fetchQuery_index) begin
        _T_257_67_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_67_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h43 == io_fetchQuery_index) begin
        _T_257_67_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_68_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h44 == io_fetchQuery_index) begin
        _T_257_68_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_68_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h44 == io_fetchQuery_index) begin
        _T_257_68_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_68_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h44 == io_fetchQuery_index) begin
        _T_257_68_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_68_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h44 == io_fetchQuery_index) begin
        _T_257_68_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_69_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h45 == io_fetchQuery_index) begin
        _T_257_69_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_69_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h45 == io_fetchQuery_index) begin
        _T_257_69_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_69_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h45 == io_fetchQuery_index) begin
        _T_257_69_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_69_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h45 == io_fetchQuery_index) begin
        _T_257_69_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_70_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h46 == io_fetchQuery_index) begin
        _T_257_70_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_70_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h46 == io_fetchQuery_index) begin
        _T_257_70_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_70_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h46 == io_fetchQuery_index) begin
        _T_257_70_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_70_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h46 == io_fetchQuery_index) begin
        _T_257_70_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_71_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h47 == io_fetchQuery_index) begin
        _T_257_71_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_71_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h47 == io_fetchQuery_index) begin
        _T_257_71_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_71_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h47 == io_fetchQuery_index) begin
        _T_257_71_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_71_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h47 == io_fetchQuery_index) begin
        _T_257_71_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_72_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h48 == io_fetchQuery_index) begin
        _T_257_72_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_72_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h48 == io_fetchQuery_index) begin
        _T_257_72_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_72_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h48 == io_fetchQuery_index) begin
        _T_257_72_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_72_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h48 == io_fetchQuery_index) begin
        _T_257_72_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_73_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h49 == io_fetchQuery_index) begin
        _T_257_73_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_73_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h49 == io_fetchQuery_index) begin
        _T_257_73_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_73_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h49 == io_fetchQuery_index) begin
        _T_257_73_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_73_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h49 == io_fetchQuery_index) begin
        _T_257_73_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_74_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h4a == io_fetchQuery_index) begin
        _T_257_74_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_74_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h4a == io_fetchQuery_index) begin
        _T_257_74_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_74_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h4a == io_fetchQuery_index) begin
        _T_257_74_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_74_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h4a == io_fetchQuery_index) begin
        _T_257_74_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_75_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h4b == io_fetchQuery_index) begin
        _T_257_75_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_75_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h4b == io_fetchQuery_index) begin
        _T_257_75_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_75_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h4b == io_fetchQuery_index) begin
        _T_257_75_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_75_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h4b == io_fetchQuery_index) begin
        _T_257_75_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_76_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h4c == io_fetchQuery_index) begin
        _T_257_76_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_76_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h4c == io_fetchQuery_index) begin
        _T_257_76_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_76_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h4c == io_fetchQuery_index) begin
        _T_257_76_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_76_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h4c == io_fetchQuery_index) begin
        _T_257_76_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_77_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h4d == io_fetchQuery_index) begin
        _T_257_77_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_77_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h4d == io_fetchQuery_index) begin
        _T_257_77_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_77_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h4d == io_fetchQuery_index) begin
        _T_257_77_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_77_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h4d == io_fetchQuery_index) begin
        _T_257_77_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_78_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h4e == io_fetchQuery_index) begin
        _T_257_78_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_78_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h4e == io_fetchQuery_index) begin
        _T_257_78_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_78_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h4e == io_fetchQuery_index) begin
        _T_257_78_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_78_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h4e == io_fetchQuery_index) begin
        _T_257_78_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_79_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h4f == io_fetchQuery_index) begin
        _T_257_79_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_79_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h4f == io_fetchQuery_index) begin
        _T_257_79_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_79_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h4f == io_fetchQuery_index) begin
        _T_257_79_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_79_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h4f == io_fetchQuery_index) begin
        _T_257_79_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_80_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h50 == io_fetchQuery_index) begin
        _T_257_80_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_80_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h50 == io_fetchQuery_index) begin
        _T_257_80_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_80_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h50 == io_fetchQuery_index) begin
        _T_257_80_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_80_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h50 == io_fetchQuery_index) begin
        _T_257_80_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_81_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h51 == io_fetchQuery_index) begin
        _T_257_81_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_81_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h51 == io_fetchQuery_index) begin
        _T_257_81_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_81_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h51 == io_fetchQuery_index) begin
        _T_257_81_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_81_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h51 == io_fetchQuery_index) begin
        _T_257_81_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_82_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h52 == io_fetchQuery_index) begin
        _T_257_82_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_82_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h52 == io_fetchQuery_index) begin
        _T_257_82_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_82_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h52 == io_fetchQuery_index) begin
        _T_257_82_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_82_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h52 == io_fetchQuery_index) begin
        _T_257_82_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_83_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h53 == io_fetchQuery_index) begin
        _T_257_83_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_83_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h53 == io_fetchQuery_index) begin
        _T_257_83_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_83_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h53 == io_fetchQuery_index) begin
        _T_257_83_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_83_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h53 == io_fetchQuery_index) begin
        _T_257_83_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_84_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h54 == io_fetchQuery_index) begin
        _T_257_84_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_84_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h54 == io_fetchQuery_index) begin
        _T_257_84_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_84_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h54 == io_fetchQuery_index) begin
        _T_257_84_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_84_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h54 == io_fetchQuery_index) begin
        _T_257_84_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_85_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h55 == io_fetchQuery_index) begin
        _T_257_85_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_85_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h55 == io_fetchQuery_index) begin
        _T_257_85_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_85_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h55 == io_fetchQuery_index) begin
        _T_257_85_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_85_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h55 == io_fetchQuery_index) begin
        _T_257_85_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_86_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h56 == io_fetchQuery_index) begin
        _T_257_86_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_86_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h56 == io_fetchQuery_index) begin
        _T_257_86_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_86_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h56 == io_fetchQuery_index) begin
        _T_257_86_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_86_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h56 == io_fetchQuery_index) begin
        _T_257_86_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_87_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h57 == io_fetchQuery_index) begin
        _T_257_87_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_87_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h57 == io_fetchQuery_index) begin
        _T_257_87_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_87_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h57 == io_fetchQuery_index) begin
        _T_257_87_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_87_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h57 == io_fetchQuery_index) begin
        _T_257_87_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_88_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h58 == io_fetchQuery_index) begin
        _T_257_88_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_88_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h58 == io_fetchQuery_index) begin
        _T_257_88_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_88_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h58 == io_fetchQuery_index) begin
        _T_257_88_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_88_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h58 == io_fetchQuery_index) begin
        _T_257_88_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_89_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h59 == io_fetchQuery_index) begin
        _T_257_89_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_89_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h59 == io_fetchQuery_index) begin
        _T_257_89_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_89_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h59 == io_fetchQuery_index) begin
        _T_257_89_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_89_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h59 == io_fetchQuery_index) begin
        _T_257_89_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_90_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h5a == io_fetchQuery_index) begin
        _T_257_90_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_90_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h5a == io_fetchQuery_index) begin
        _T_257_90_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_90_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h5a == io_fetchQuery_index) begin
        _T_257_90_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_90_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h5a == io_fetchQuery_index) begin
        _T_257_90_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_91_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h5b == io_fetchQuery_index) begin
        _T_257_91_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_91_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h5b == io_fetchQuery_index) begin
        _T_257_91_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_91_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h5b == io_fetchQuery_index) begin
        _T_257_91_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_91_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h5b == io_fetchQuery_index) begin
        _T_257_91_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_92_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h5c == io_fetchQuery_index) begin
        _T_257_92_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_92_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h5c == io_fetchQuery_index) begin
        _T_257_92_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_92_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h5c == io_fetchQuery_index) begin
        _T_257_92_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_92_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h5c == io_fetchQuery_index) begin
        _T_257_92_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_93_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h5d == io_fetchQuery_index) begin
        _T_257_93_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_93_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h5d == io_fetchQuery_index) begin
        _T_257_93_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_93_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h5d == io_fetchQuery_index) begin
        _T_257_93_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_93_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h5d == io_fetchQuery_index) begin
        _T_257_93_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_94_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h5e == io_fetchQuery_index) begin
        _T_257_94_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_94_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h5e == io_fetchQuery_index) begin
        _T_257_94_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_94_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h5e == io_fetchQuery_index) begin
        _T_257_94_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_94_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h5e == io_fetchQuery_index) begin
        _T_257_94_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_95_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h5f == io_fetchQuery_index) begin
        _T_257_95_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_95_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h5f == io_fetchQuery_index) begin
        _T_257_95_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_95_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h5f == io_fetchQuery_index) begin
        _T_257_95_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_95_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h5f == io_fetchQuery_index) begin
        _T_257_95_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_96_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h60 == io_fetchQuery_index) begin
        _T_257_96_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_96_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h60 == io_fetchQuery_index) begin
        _T_257_96_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_96_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h60 == io_fetchQuery_index) begin
        _T_257_96_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_96_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h60 == io_fetchQuery_index) begin
        _T_257_96_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_97_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h61 == io_fetchQuery_index) begin
        _T_257_97_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_97_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h61 == io_fetchQuery_index) begin
        _T_257_97_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_97_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h61 == io_fetchQuery_index) begin
        _T_257_97_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_97_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h61 == io_fetchQuery_index) begin
        _T_257_97_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_98_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h62 == io_fetchQuery_index) begin
        _T_257_98_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_98_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h62 == io_fetchQuery_index) begin
        _T_257_98_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_98_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h62 == io_fetchQuery_index) begin
        _T_257_98_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_98_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h62 == io_fetchQuery_index) begin
        _T_257_98_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_99_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h63 == io_fetchQuery_index) begin
        _T_257_99_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_99_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h63 == io_fetchQuery_index) begin
        _T_257_99_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_99_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h63 == io_fetchQuery_index) begin
        _T_257_99_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_99_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h63 == io_fetchQuery_index) begin
        _T_257_99_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_100_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h64 == io_fetchQuery_index) begin
        _T_257_100_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_100_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h64 == io_fetchQuery_index) begin
        _T_257_100_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_100_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h64 == io_fetchQuery_index) begin
        _T_257_100_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_100_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h64 == io_fetchQuery_index) begin
        _T_257_100_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_101_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h65 == io_fetchQuery_index) begin
        _T_257_101_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_101_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h65 == io_fetchQuery_index) begin
        _T_257_101_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_101_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h65 == io_fetchQuery_index) begin
        _T_257_101_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_101_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h65 == io_fetchQuery_index) begin
        _T_257_101_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_102_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h66 == io_fetchQuery_index) begin
        _T_257_102_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_102_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h66 == io_fetchQuery_index) begin
        _T_257_102_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_102_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h66 == io_fetchQuery_index) begin
        _T_257_102_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_102_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h66 == io_fetchQuery_index) begin
        _T_257_102_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_103_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h67 == io_fetchQuery_index) begin
        _T_257_103_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_103_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h67 == io_fetchQuery_index) begin
        _T_257_103_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_103_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h67 == io_fetchQuery_index) begin
        _T_257_103_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_103_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h67 == io_fetchQuery_index) begin
        _T_257_103_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_104_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h68 == io_fetchQuery_index) begin
        _T_257_104_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_104_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h68 == io_fetchQuery_index) begin
        _T_257_104_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_104_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h68 == io_fetchQuery_index) begin
        _T_257_104_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_104_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h68 == io_fetchQuery_index) begin
        _T_257_104_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_105_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h69 == io_fetchQuery_index) begin
        _T_257_105_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_105_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h69 == io_fetchQuery_index) begin
        _T_257_105_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_105_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h69 == io_fetchQuery_index) begin
        _T_257_105_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_105_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h69 == io_fetchQuery_index) begin
        _T_257_105_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_106_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h6a == io_fetchQuery_index) begin
        _T_257_106_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_106_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h6a == io_fetchQuery_index) begin
        _T_257_106_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_106_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h6a == io_fetchQuery_index) begin
        _T_257_106_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_106_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h6a == io_fetchQuery_index) begin
        _T_257_106_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_107_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h6b == io_fetchQuery_index) begin
        _T_257_107_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_107_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h6b == io_fetchQuery_index) begin
        _T_257_107_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_107_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h6b == io_fetchQuery_index) begin
        _T_257_107_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_107_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h6b == io_fetchQuery_index) begin
        _T_257_107_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_108_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h6c == io_fetchQuery_index) begin
        _T_257_108_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_108_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h6c == io_fetchQuery_index) begin
        _T_257_108_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_108_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h6c == io_fetchQuery_index) begin
        _T_257_108_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_108_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h6c == io_fetchQuery_index) begin
        _T_257_108_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_109_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h6d == io_fetchQuery_index) begin
        _T_257_109_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_109_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h6d == io_fetchQuery_index) begin
        _T_257_109_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_109_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h6d == io_fetchQuery_index) begin
        _T_257_109_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_109_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h6d == io_fetchQuery_index) begin
        _T_257_109_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_110_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h6e == io_fetchQuery_index) begin
        _T_257_110_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_110_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h6e == io_fetchQuery_index) begin
        _T_257_110_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_110_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h6e == io_fetchQuery_index) begin
        _T_257_110_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_110_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h6e == io_fetchQuery_index) begin
        _T_257_110_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_111_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h6f == io_fetchQuery_index) begin
        _T_257_111_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_111_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h6f == io_fetchQuery_index) begin
        _T_257_111_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_111_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h6f == io_fetchQuery_index) begin
        _T_257_111_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_111_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h6f == io_fetchQuery_index) begin
        _T_257_111_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_112_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h70 == io_fetchQuery_index) begin
        _T_257_112_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_112_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h70 == io_fetchQuery_index) begin
        _T_257_112_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_112_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h70 == io_fetchQuery_index) begin
        _T_257_112_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_112_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h70 == io_fetchQuery_index) begin
        _T_257_112_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_113_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h71 == io_fetchQuery_index) begin
        _T_257_113_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_113_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h71 == io_fetchQuery_index) begin
        _T_257_113_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_113_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h71 == io_fetchQuery_index) begin
        _T_257_113_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_113_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h71 == io_fetchQuery_index) begin
        _T_257_113_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_114_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h72 == io_fetchQuery_index) begin
        _T_257_114_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_114_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h72 == io_fetchQuery_index) begin
        _T_257_114_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_114_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h72 == io_fetchQuery_index) begin
        _T_257_114_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_114_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h72 == io_fetchQuery_index) begin
        _T_257_114_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_115_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h73 == io_fetchQuery_index) begin
        _T_257_115_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_115_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h73 == io_fetchQuery_index) begin
        _T_257_115_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_115_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h73 == io_fetchQuery_index) begin
        _T_257_115_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_115_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h73 == io_fetchQuery_index) begin
        _T_257_115_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_116_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h74 == io_fetchQuery_index) begin
        _T_257_116_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_116_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h74 == io_fetchQuery_index) begin
        _T_257_116_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_116_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h74 == io_fetchQuery_index) begin
        _T_257_116_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_116_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h74 == io_fetchQuery_index) begin
        _T_257_116_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_117_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h75 == io_fetchQuery_index) begin
        _T_257_117_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_117_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h75 == io_fetchQuery_index) begin
        _T_257_117_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_117_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h75 == io_fetchQuery_index) begin
        _T_257_117_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_117_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h75 == io_fetchQuery_index) begin
        _T_257_117_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_118_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h76 == io_fetchQuery_index) begin
        _T_257_118_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_118_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h76 == io_fetchQuery_index) begin
        _T_257_118_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_118_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h76 == io_fetchQuery_index) begin
        _T_257_118_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_118_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h76 == io_fetchQuery_index) begin
        _T_257_118_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_119_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h77 == io_fetchQuery_index) begin
        _T_257_119_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_119_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h77 == io_fetchQuery_index) begin
        _T_257_119_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_119_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h77 == io_fetchQuery_index) begin
        _T_257_119_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_119_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h77 == io_fetchQuery_index) begin
        _T_257_119_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_120_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h78 == io_fetchQuery_index) begin
        _T_257_120_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_120_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h78 == io_fetchQuery_index) begin
        _T_257_120_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_120_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h78 == io_fetchQuery_index) begin
        _T_257_120_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_120_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h78 == io_fetchQuery_index) begin
        _T_257_120_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_121_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h79 == io_fetchQuery_index) begin
        _T_257_121_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_121_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h79 == io_fetchQuery_index) begin
        _T_257_121_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_121_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h79 == io_fetchQuery_index) begin
        _T_257_121_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_121_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h79 == io_fetchQuery_index) begin
        _T_257_121_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_122_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h7a == io_fetchQuery_index) begin
        _T_257_122_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_122_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h7a == io_fetchQuery_index) begin
        _T_257_122_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_122_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h7a == io_fetchQuery_index) begin
        _T_257_122_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_122_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h7a == io_fetchQuery_index) begin
        _T_257_122_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_123_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h7b == io_fetchQuery_index) begin
        _T_257_123_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_123_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h7b == io_fetchQuery_index) begin
        _T_257_123_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_123_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h7b == io_fetchQuery_index) begin
        _T_257_123_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_123_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h7b == io_fetchQuery_index) begin
        _T_257_123_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_124_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h7c == io_fetchQuery_index) begin
        _T_257_124_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_124_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h7c == io_fetchQuery_index) begin
        _T_257_124_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_124_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h7c == io_fetchQuery_index) begin
        _T_257_124_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_124_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h7c == io_fetchQuery_index) begin
        _T_257_124_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_125_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h7d == io_fetchQuery_index) begin
        _T_257_125_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_125_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h7d == io_fetchQuery_index) begin
        _T_257_125_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_125_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h7d == io_fetchQuery_index) begin
        _T_257_125_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_125_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h7d == io_fetchQuery_index) begin
        _T_257_125_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_126_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h7e == io_fetchQuery_index) begin
        _T_257_126_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_126_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h7e == io_fetchQuery_index) begin
        _T_257_126_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_126_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h7e == io_fetchQuery_index) begin
        _T_257_126_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_126_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h7e == io_fetchQuery_index) begin
        _T_257_126_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_127_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h7f == io_fetchQuery_index) begin
        _T_257_127_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_127_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h7f == io_fetchQuery_index) begin
        _T_257_127_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_127_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h7f == io_fetchQuery_index) begin
        _T_257_127_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_127_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h7f == io_fetchQuery_index) begin
        _T_257_127_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_128_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h80 == io_fetchQuery_index) begin
        _T_257_128_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_128_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h80 == io_fetchQuery_index) begin
        _T_257_128_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_128_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h80 == io_fetchQuery_index) begin
        _T_257_128_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_128_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h80 == io_fetchQuery_index) begin
        _T_257_128_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_129_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h81 == io_fetchQuery_index) begin
        _T_257_129_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_129_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h81 == io_fetchQuery_index) begin
        _T_257_129_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_129_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h81 == io_fetchQuery_index) begin
        _T_257_129_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_129_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h81 == io_fetchQuery_index) begin
        _T_257_129_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_130_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h82 == io_fetchQuery_index) begin
        _T_257_130_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_130_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h82 == io_fetchQuery_index) begin
        _T_257_130_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_130_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h82 == io_fetchQuery_index) begin
        _T_257_130_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_130_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h82 == io_fetchQuery_index) begin
        _T_257_130_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_131_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h83 == io_fetchQuery_index) begin
        _T_257_131_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_131_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h83 == io_fetchQuery_index) begin
        _T_257_131_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_131_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h83 == io_fetchQuery_index) begin
        _T_257_131_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_131_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h83 == io_fetchQuery_index) begin
        _T_257_131_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_132_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h84 == io_fetchQuery_index) begin
        _T_257_132_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_132_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h84 == io_fetchQuery_index) begin
        _T_257_132_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_132_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h84 == io_fetchQuery_index) begin
        _T_257_132_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_132_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h84 == io_fetchQuery_index) begin
        _T_257_132_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_133_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h85 == io_fetchQuery_index) begin
        _T_257_133_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_133_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h85 == io_fetchQuery_index) begin
        _T_257_133_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_133_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h85 == io_fetchQuery_index) begin
        _T_257_133_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_133_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h85 == io_fetchQuery_index) begin
        _T_257_133_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_134_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h86 == io_fetchQuery_index) begin
        _T_257_134_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_134_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h86 == io_fetchQuery_index) begin
        _T_257_134_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_134_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h86 == io_fetchQuery_index) begin
        _T_257_134_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_134_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h86 == io_fetchQuery_index) begin
        _T_257_134_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_135_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h87 == io_fetchQuery_index) begin
        _T_257_135_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_135_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h87 == io_fetchQuery_index) begin
        _T_257_135_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_135_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h87 == io_fetchQuery_index) begin
        _T_257_135_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_135_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h87 == io_fetchQuery_index) begin
        _T_257_135_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_136_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h88 == io_fetchQuery_index) begin
        _T_257_136_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_136_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h88 == io_fetchQuery_index) begin
        _T_257_136_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_136_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h88 == io_fetchQuery_index) begin
        _T_257_136_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_136_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h88 == io_fetchQuery_index) begin
        _T_257_136_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_137_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h89 == io_fetchQuery_index) begin
        _T_257_137_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_137_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h89 == io_fetchQuery_index) begin
        _T_257_137_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_137_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h89 == io_fetchQuery_index) begin
        _T_257_137_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_137_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h89 == io_fetchQuery_index) begin
        _T_257_137_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_138_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h8a == io_fetchQuery_index) begin
        _T_257_138_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_138_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h8a == io_fetchQuery_index) begin
        _T_257_138_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_138_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h8a == io_fetchQuery_index) begin
        _T_257_138_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_138_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h8a == io_fetchQuery_index) begin
        _T_257_138_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_139_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h8b == io_fetchQuery_index) begin
        _T_257_139_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_139_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h8b == io_fetchQuery_index) begin
        _T_257_139_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_139_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h8b == io_fetchQuery_index) begin
        _T_257_139_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_139_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h8b == io_fetchQuery_index) begin
        _T_257_139_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_140_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h8c == io_fetchQuery_index) begin
        _T_257_140_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_140_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h8c == io_fetchQuery_index) begin
        _T_257_140_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_140_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h8c == io_fetchQuery_index) begin
        _T_257_140_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_140_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h8c == io_fetchQuery_index) begin
        _T_257_140_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_141_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h8d == io_fetchQuery_index) begin
        _T_257_141_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_141_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h8d == io_fetchQuery_index) begin
        _T_257_141_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_141_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h8d == io_fetchQuery_index) begin
        _T_257_141_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_141_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h8d == io_fetchQuery_index) begin
        _T_257_141_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_142_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h8e == io_fetchQuery_index) begin
        _T_257_142_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_142_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h8e == io_fetchQuery_index) begin
        _T_257_142_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_142_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h8e == io_fetchQuery_index) begin
        _T_257_142_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_142_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h8e == io_fetchQuery_index) begin
        _T_257_142_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_143_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h8f == io_fetchQuery_index) begin
        _T_257_143_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_143_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h8f == io_fetchQuery_index) begin
        _T_257_143_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_143_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h8f == io_fetchQuery_index) begin
        _T_257_143_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_143_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h8f == io_fetchQuery_index) begin
        _T_257_143_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_144_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h90 == io_fetchQuery_index) begin
        _T_257_144_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_144_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h90 == io_fetchQuery_index) begin
        _T_257_144_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_144_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h90 == io_fetchQuery_index) begin
        _T_257_144_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_144_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h90 == io_fetchQuery_index) begin
        _T_257_144_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_145_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h91 == io_fetchQuery_index) begin
        _T_257_145_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_145_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h91 == io_fetchQuery_index) begin
        _T_257_145_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_145_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h91 == io_fetchQuery_index) begin
        _T_257_145_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_145_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h91 == io_fetchQuery_index) begin
        _T_257_145_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_146_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h92 == io_fetchQuery_index) begin
        _T_257_146_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_146_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h92 == io_fetchQuery_index) begin
        _T_257_146_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_146_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h92 == io_fetchQuery_index) begin
        _T_257_146_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_146_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h92 == io_fetchQuery_index) begin
        _T_257_146_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_147_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h93 == io_fetchQuery_index) begin
        _T_257_147_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_147_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h93 == io_fetchQuery_index) begin
        _T_257_147_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_147_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h93 == io_fetchQuery_index) begin
        _T_257_147_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_147_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h93 == io_fetchQuery_index) begin
        _T_257_147_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_148_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h94 == io_fetchQuery_index) begin
        _T_257_148_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_148_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h94 == io_fetchQuery_index) begin
        _T_257_148_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_148_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h94 == io_fetchQuery_index) begin
        _T_257_148_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_148_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h94 == io_fetchQuery_index) begin
        _T_257_148_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_149_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h95 == io_fetchQuery_index) begin
        _T_257_149_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_149_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h95 == io_fetchQuery_index) begin
        _T_257_149_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_149_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h95 == io_fetchQuery_index) begin
        _T_257_149_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_149_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h95 == io_fetchQuery_index) begin
        _T_257_149_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_150_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h96 == io_fetchQuery_index) begin
        _T_257_150_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_150_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h96 == io_fetchQuery_index) begin
        _T_257_150_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_150_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h96 == io_fetchQuery_index) begin
        _T_257_150_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_150_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h96 == io_fetchQuery_index) begin
        _T_257_150_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_151_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h97 == io_fetchQuery_index) begin
        _T_257_151_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_151_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h97 == io_fetchQuery_index) begin
        _T_257_151_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_151_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h97 == io_fetchQuery_index) begin
        _T_257_151_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_151_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h97 == io_fetchQuery_index) begin
        _T_257_151_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_152_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h98 == io_fetchQuery_index) begin
        _T_257_152_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_152_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h98 == io_fetchQuery_index) begin
        _T_257_152_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_152_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h98 == io_fetchQuery_index) begin
        _T_257_152_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_152_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h98 == io_fetchQuery_index) begin
        _T_257_152_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_153_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h99 == io_fetchQuery_index) begin
        _T_257_153_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_153_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h99 == io_fetchQuery_index) begin
        _T_257_153_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_153_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h99 == io_fetchQuery_index) begin
        _T_257_153_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_153_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h99 == io_fetchQuery_index) begin
        _T_257_153_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_154_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h9a == io_fetchQuery_index) begin
        _T_257_154_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_154_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h9a == io_fetchQuery_index) begin
        _T_257_154_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_154_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h9a == io_fetchQuery_index) begin
        _T_257_154_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_154_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h9a == io_fetchQuery_index) begin
        _T_257_154_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_155_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h9b == io_fetchQuery_index) begin
        _T_257_155_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_155_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h9b == io_fetchQuery_index) begin
        _T_257_155_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_155_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h9b == io_fetchQuery_index) begin
        _T_257_155_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_155_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h9b == io_fetchQuery_index) begin
        _T_257_155_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_156_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h9c == io_fetchQuery_index) begin
        _T_257_156_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_156_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h9c == io_fetchQuery_index) begin
        _T_257_156_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_156_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h9c == io_fetchQuery_index) begin
        _T_257_156_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_156_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h9c == io_fetchQuery_index) begin
        _T_257_156_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_157_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h9d == io_fetchQuery_index) begin
        _T_257_157_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_157_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h9d == io_fetchQuery_index) begin
        _T_257_157_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_157_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h9d == io_fetchQuery_index) begin
        _T_257_157_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_157_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h9d == io_fetchQuery_index) begin
        _T_257_157_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_158_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h9e == io_fetchQuery_index) begin
        _T_257_158_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_158_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h9e == io_fetchQuery_index) begin
        _T_257_158_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_158_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h9e == io_fetchQuery_index) begin
        _T_257_158_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_158_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h9e == io_fetchQuery_index) begin
        _T_257_158_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_159_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h9f == io_fetchQuery_index) begin
        _T_257_159_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_159_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h9f == io_fetchQuery_index) begin
        _T_257_159_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_159_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h9f == io_fetchQuery_index) begin
        _T_257_159_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_159_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'h9f == io_fetchQuery_index) begin
        _T_257_159_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_160_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'ha0 == io_fetchQuery_index) begin
        _T_257_160_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_160_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'ha0 == io_fetchQuery_index) begin
        _T_257_160_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_160_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'ha0 == io_fetchQuery_index) begin
        _T_257_160_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_160_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'ha0 == io_fetchQuery_index) begin
        _T_257_160_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_161_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'ha1 == io_fetchQuery_index) begin
        _T_257_161_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_161_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'ha1 == io_fetchQuery_index) begin
        _T_257_161_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_161_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'ha1 == io_fetchQuery_index) begin
        _T_257_161_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_161_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'ha1 == io_fetchQuery_index) begin
        _T_257_161_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_162_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'ha2 == io_fetchQuery_index) begin
        _T_257_162_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_162_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'ha2 == io_fetchQuery_index) begin
        _T_257_162_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_162_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'ha2 == io_fetchQuery_index) begin
        _T_257_162_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_162_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'ha2 == io_fetchQuery_index) begin
        _T_257_162_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_163_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'ha3 == io_fetchQuery_index) begin
        _T_257_163_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_163_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'ha3 == io_fetchQuery_index) begin
        _T_257_163_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_163_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'ha3 == io_fetchQuery_index) begin
        _T_257_163_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_163_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'ha3 == io_fetchQuery_index) begin
        _T_257_163_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_164_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'ha4 == io_fetchQuery_index) begin
        _T_257_164_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_164_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'ha4 == io_fetchQuery_index) begin
        _T_257_164_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_164_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'ha4 == io_fetchQuery_index) begin
        _T_257_164_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_164_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'ha4 == io_fetchQuery_index) begin
        _T_257_164_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_165_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'ha5 == io_fetchQuery_index) begin
        _T_257_165_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_165_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'ha5 == io_fetchQuery_index) begin
        _T_257_165_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_165_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'ha5 == io_fetchQuery_index) begin
        _T_257_165_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_165_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'ha5 == io_fetchQuery_index) begin
        _T_257_165_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_166_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'ha6 == io_fetchQuery_index) begin
        _T_257_166_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_166_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'ha6 == io_fetchQuery_index) begin
        _T_257_166_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_166_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'ha6 == io_fetchQuery_index) begin
        _T_257_166_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_166_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'ha6 == io_fetchQuery_index) begin
        _T_257_166_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_167_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'ha7 == io_fetchQuery_index) begin
        _T_257_167_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_167_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'ha7 == io_fetchQuery_index) begin
        _T_257_167_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_167_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'ha7 == io_fetchQuery_index) begin
        _T_257_167_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_167_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'ha7 == io_fetchQuery_index) begin
        _T_257_167_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_168_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'ha8 == io_fetchQuery_index) begin
        _T_257_168_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_168_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'ha8 == io_fetchQuery_index) begin
        _T_257_168_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_168_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'ha8 == io_fetchQuery_index) begin
        _T_257_168_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_168_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'ha8 == io_fetchQuery_index) begin
        _T_257_168_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_169_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'ha9 == io_fetchQuery_index) begin
        _T_257_169_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_169_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'ha9 == io_fetchQuery_index) begin
        _T_257_169_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_169_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'ha9 == io_fetchQuery_index) begin
        _T_257_169_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_169_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'ha9 == io_fetchQuery_index) begin
        _T_257_169_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_170_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'haa == io_fetchQuery_index) begin
        _T_257_170_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_170_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'haa == io_fetchQuery_index) begin
        _T_257_170_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_170_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'haa == io_fetchQuery_index) begin
        _T_257_170_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_170_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'haa == io_fetchQuery_index) begin
        _T_257_170_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_171_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hab == io_fetchQuery_index) begin
        _T_257_171_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_171_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hab == io_fetchQuery_index) begin
        _T_257_171_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_171_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hab == io_fetchQuery_index) begin
        _T_257_171_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_171_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hab == io_fetchQuery_index) begin
        _T_257_171_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_172_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hac == io_fetchQuery_index) begin
        _T_257_172_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_172_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hac == io_fetchQuery_index) begin
        _T_257_172_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_172_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hac == io_fetchQuery_index) begin
        _T_257_172_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_172_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hac == io_fetchQuery_index) begin
        _T_257_172_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_173_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'had == io_fetchQuery_index) begin
        _T_257_173_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_173_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'had == io_fetchQuery_index) begin
        _T_257_173_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_173_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'had == io_fetchQuery_index) begin
        _T_257_173_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_173_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'had == io_fetchQuery_index) begin
        _T_257_173_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_174_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hae == io_fetchQuery_index) begin
        _T_257_174_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_174_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hae == io_fetchQuery_index) begin
        _T_257_174_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_174_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hae == io_fetchQuery_index) begin
        _T_257_174_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_174_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hae == io_fetchQuery_index) begin
        _T_257_174_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_175_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'haf == io_fetchQuery_index) begin
        _T_257_175_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_175_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'haf == io_fetchQuery_index) begin
        _T_257_175_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_175_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'haf == io_fetchQuery_index) begin
        _T_257_175_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_175_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'haf == io_fetchQuery_index) begin
        _T_257_175_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_176_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hb0 == io_fetchQuery_index) begin
        _T_257_176_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_176_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hb0 == io_fetchQuery_index) begin
        _T_257_176_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_176_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hb0 == io_fetchQuery_index) begin
        _T_257_176_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_176_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hb0 == io_fetchQuery_index) begin
        _T_257_176_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_177_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hb1 == io_fetchQuery_index) begin
        _T_257_177_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_177_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hb1 == io_fetchQuery_index) begin
        _T_257_177_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_177_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hb1 == io_fetchQuery_index) begin
        _T_257_177_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_177_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hb1 == io_fetchQuery_index) begin
        _T_257_177_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_178_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hb2 == io_fetchQuery_index) begin
        _T_257_178_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_178_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hb2 == io_fetchQuery_index) begin
        _T_257_178_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_178_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hb2 == io_fetchQuery_index) begin
        _T_257_178_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_178_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hb2 == io_fetchQuery_index) begin
        _T_257_178_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_179_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hb3 == io_fetchQuery_index) begin
        _T_257_179_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_179_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hb3 == io_fetchQuery_index) begin
        _T_257_179_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_179_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hb3 == io_fetchQuery_index) begin
        _T_257_179_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_179_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hb3 == io_fetchQuery_index) begin
        _T_257_179_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_180_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hb4 == io_fetchQuery_index) begin
        _T_257_180_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_180_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hb4 == io_fetchQuery_index) begin
        _T_257_180_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_180_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hb4 == io_fetchQuery_index) begin
        _T_257_180_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_180_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hb4 == io_fetchQuery_index) begin
        _T_257_180_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_181_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hb5 == io_fetchQuery_index) begin
        _T_257_181_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_181_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hb5 == io_fetchQuery_index) begin
        _T_257_181_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_181_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hb5 == io_fetchQuery_index) begin
        _T_257_181_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_181_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hb5 == io_fetchQuery_index) begin
        _T_257_181_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_182_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hb6 == io_fetchQuery_index) begin
        _T_257_182_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_182_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hb6 == io_fetchQuery_index) begin
        _T_257_182_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_182_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hb6 == io_fetchQuery_index) begin
        _T_257_182_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_182_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hb6 == io_fetchQuery_index) begin
        _T_257_182_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_183_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hb7 == io_fetchQuery_index) begin
        _T_257_183_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_183_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hb7 == io_fetchQuery_index) begin
        _T_257_183_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_183_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hb7 == io_fetchQuery_index) begin
        _T_257_183_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_183_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hb7 == io_fetchQuery_index) begin
        _T_257_183_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_184_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hb8 == io_fetchQuery_index) begin
        _T_257_184_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_184_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hb8 == io_fetchQuery_index) begin
        _T_257_184_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_184_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hb8 == io_fetchQuery_index) begin
        _T_257_184_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_184_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hb8 == io_fetchQuery_index) begin
        _T_257_184_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_185_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hb9 == io_fetchQuery_index) begin
        _T_257_185_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_185_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hb9 == io_fetchQuery_index) begin
        _T_257_185_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_185_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hb9 == io_fetchQuery_index) begin
        _T_257_185_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_185_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hb9 == io_fetchQuery_index) begin
        _T_257_185_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_186_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hba == io_fetchQuery_index) begin
        _T_257_186_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_186_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hba == io_fetchQuery_index) begin
        _T_257_186_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_186_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hba == io_fetchQuery_index) begin
        _T_257_186_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_186_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hba == io_fetchQuery_index) begin
        _T_257_186_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_187_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hbb == io_fetchQuery_index) begin
        _T_257_187_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_187_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hbb == io_fetchQuery_index) begin
        _T_257_187_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_187_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hbb == io_fetchQuery_index) begin
        _T_257_187_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_187_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hbb == io_fetchQuery_index) begin
        _T_257_187_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_188_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hbc == io_fetchQuery_index) begin
        _T_257_188_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_188_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hbc == io_fetchQuery_index) begin
        _T_257_188_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_188_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hbc == io_fetchQuery_index) begin
        _T_257_188_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_188_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hbc == io_fetchQuery_index) begin
        _T_257_188_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_189_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hbd == io_fetchQuery_index) begin
        _T_257_189_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_189_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hbd == io_fetchQuery_index) begin
        _T_257_189_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_189_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hbd == io_fetchQuery_index) begin
        _T_257_189_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_189_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hbd == io_fetchQuery_index) begin
        _T_257_189_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_190_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hbe == io_fetchQuery_index) begin
        _T_257_190_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_190_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hbe == io_fetchQuery_index) begin
        _T_257_190_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_190_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hbe == io_fetchQuery_index) begin
        _T_257_190_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_190_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hbe == io_fetchQuery_index) begin
        _T_257_190_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_191_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hbf == io_fetchQuery_index) begin
        _T_257_191_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_191_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hbf == io_fetchQuery_index) begin
        _T_257_191_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_191_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hbf == io_fetchQuery_index) begin
        _T_257_191_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_191_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hbf == io_fetchQuery_index) begin
        _T_257_191_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_192_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hc0 == io_fetchQuery_index) begin
        _T_257_192_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_192_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hc0 == io_fetchQuery_index) begin
        _T_257_192_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_192_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hc0 == io_fetchQuery_index) begin
        _T_257_192_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_192_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hc0 == io_fetchQuery_index) begin
        _T_257_192_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_193_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hc1 == io_fetchQuery_index) begin
        _T_257_193_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_193_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hc1 == io_fetchQuery_index) begin
        _T_257_193_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_193_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hc1 == io_fetchQuery_index) begin
        _T_257_193_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_193_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hc1 == io_fetchQuery_index) begin
        _T_257_193_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_194_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hc2 == io_fetchQuery_index) begin
        _T_257_194_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_194_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hc2 == io_fetchQuery_index) begin
        _T_257_194_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_194_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hc2 == io_fetchQuery_index) begin
        _T_257_194_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_194_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hc2 == io_fetchQuery_index) begin
        _T_257_194_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_195_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hc3 == io_fetchQuery_index) begin
        _T_257_195_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_195_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hc3 == io_fetchQuery_index) begin
        _T_257_195_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_195_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hc3 == io_fetchQuery_index) begin
        _T_257_195_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_195_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hc3 == io_fetchQuery_index) begin
        _T_257_195_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_196_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hc4 == io_fetchQuery_index) begin
        _T_257_196_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_196_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hc4 == io_fetchQuery_index) begin
        _T_257_196_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_196_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hc4 == io_fetchQuery_index) begin
        _T_257_196_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_196_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hc4 == io_fetchQuery_index) begin
        _T_257_196_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_197_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hc5 == io_fetchQuery_index) begin
        _T_257_197_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_197_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hc5 == io_fetchQuery_index) begin
        _T_257_197_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_197_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hc5 == io_fetchQuery_index) begin
        _T_257_197_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_197_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hc5 == io_fetchQuery_index) begin
        _T_257_197_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_198_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hc6 == io_fetchQuery_index) begin
        _T_257_198_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_198_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hc6 == io_fetchQuery_index) begin
        _T_257_198_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_198_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hc6 == io_fetchQuery_index) begin
        _T_257_198_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_198_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hc6 == io_fetchQuery_index) begin
        _T_257_198_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_199_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hc7 == io_fetchQuery_index) begin
        _T_257_199_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_199_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hc7 == io_fetchQuery_index) begin
        _T_257_199_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_199_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hc7 == io_fetchQuery_index) begin
        _T_257_199_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_199_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hc7 == io_fetchQuery_index) begin
        _T_257_199_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_200_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hc8 == io_fetchQuery_index) begin
        _T_257_200_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_200_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hc8 == io_fetchQuery_index) begin
        _T_257_200_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_200_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hc8 == io_fetchQuery_index) begin
        _T_257_200_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_200_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hc8 == io_fetchQuery_index) begin
        _T_257_200_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_201_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hc9 == io_fetchQuery_index) begin
        _T_257_201_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_201_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hc9 == io_fetchQuery_index) begin
        _T_257_201_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_201_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hc9 == io_fetchQuery_index) begin
        _T_257_201_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_201_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hc9 == io_fetchQuery_index) begin
        _T_257_201_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_202_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hca == io_fetchQuery_index) begin
        _T_257_202_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_202_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hca == io_fetchQuery_index) begin
        _T_257_202_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_202_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hca == io_fetchQuery_index) begin
        _T_257_202_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_202_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hca == io_fetchQuery_index) begin
        _T_257_202_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_203_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hcb == io_fetchQuery_index) begin
        _T_257_203_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_203_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hcb == io_fetchQuery_index) begin
        _T_257_203_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_203_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hcb == io_fetchQuery_index) begin
        _T_257_203_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_203_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hcb == io_fetchQuery_index) begin
        _T_257_203_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_204_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hcc == io_fetchQuery_index) begin
        _T_257_204_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_204_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hcc == io_fetchQuery_index) begin
        _T_257_204_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_204_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hcc == io_fetchQuery_index) begin
        _T_257_204_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_204_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hcc == io_fetchQuery_index) begin
        _T_257_204_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_205_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hcd == io_fetchQuery_index) begin
        _T_257_205_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_205_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hcd == io_fetchQuery_index) begin
        _T_257_205_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_205_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hcd == io_fetchQuery_index) begin
        _T_257_205_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_205_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hcd == io_fetchQuery_index) begin
        _T_257_205_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_206_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hce == io_fetchQuery_index) begin
        _T_257_206_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_206_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hce == io_fetchQuery_index) begin
        _T_257_206_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_206_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hce == io_fetchQuery_index) begin
        _T_257_206_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_206_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hce == io_fetchQuery_index) begin
        _T_257_206_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_207_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hcf == io_fetchQuery_index) begin
        _T_257_207_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_207_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hcf == io_fetchQuery_index) begin
        _T_257_207_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_207_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hcf == io_fetchQuery_index) begin
        _T_257_207_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_207_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hcf == io_fetchQuery_index) begin
        _T_257_207_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_208_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hd0 == io_fetchQuery_index) begin
        _T_257_208_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_208_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hd0 == io_fetchQuery_index) begin
        _T_257_208_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_208_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hd0 == io_fetchQuery_index) begin
        _T_257_208_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_208_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hd0 == io_fetchQuery_index) begin
        _T_257_208_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_209_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hd1 == io_fetchQuery_index) begin
        _T_257_209_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_209_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hd1 == io_fetchQuery_index) begin
        _T_257_209_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_209_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hd1 == io_fetchQuery_index) begin
        _T_257_209_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_209_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hd1 == io_fetchQuery_index) begin
        _T_257_209_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_210_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hd2 == io_fetchQuery_index) begin
        _T_257_210_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_210_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hd2 == io_fetchQuery_index) begin
        _T_257_210_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_210_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hd2 == io_fetchQuery_index) begin
        _T_257_210_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_210_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hd2 == io_fetchQuery_index) begin
        _T_257_210_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_211_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hd3 == io_fetchQuery_index) begin
        _T_257_211_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_211_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hd3 == io_fetchQuery_index) begin
        _T_257_211_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_211_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hd3 == io_fetchQuery_index) begin
        _T_257_211_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_211_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hd3 == io_fetchQuery_index) begin
        _T_257_211_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_212_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hd4 == io_fetchQuery_index) begin
        _T_257_212_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_212_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hd4 == io_fetchQuery_index) begin
        _T_257_212_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_212_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hd4 == io_fetchQuery_index) begin
        _T_257_212_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_212_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hd4 == io_fetchQuery_index) begin
        _T_257_212_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_213_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hd5 == io_fetchQuery_index) begin
        _T_257_213_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_213_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hd5 == io_fetchQuery_index) begin
        _T_257_213_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_213_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hd5 == io_fetchQuery_index) begin
        _T_257_213_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_213_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hd5 == io_fetchQuery_index) begin
        _T_257_213_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_214_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hd6 == io_fetchQuery_index) begin
        _T_257_214_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_214_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hd6 == io_fetchQuery_index) begin
        _T_257_214_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_214_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hd6 == io_fetchQuery_index) begin
        _T_257_214_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_214_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hd6 == io_fetchQuery_index) begin
        _T_257_214_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_215_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hd7 == io_fetchQuery_index) begin
        _T_257_215_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_215_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hd7 == io_fetchQuery_index) begin
        _T_257_215_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_215_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hd7 == io_fetchQuery_index) begin
        _T_257_215_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_215_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hd7 == io_fetchQuery_index) begin
        _T_257_215_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_216_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hd8 == io_fetchQuery_index) begin
        _T_257_216_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_216_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hd8 == io_fetchQuery_index) begin
        _T_257_216_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_216_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hd8 == io_fetchQuery_index) begin
        _T_257_216_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_216_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hd8 == io_fetchQuery_index) begin
        _T_257_216_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_217_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hd9 == io_fetchQuery_index) begin
        _T_257_217_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_217_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hd9 == io_fetchQuery_index) begin
        _T_257_217_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_217_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hd9 == io_fetchQuery_index) begin
        _T_257_217_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_217_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hd9 == io_fetchQuery_index) begin
        _T_257_217_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_218_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hda == io_fetchQuery_index) begin
        _T_257_218_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_218_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hda == io_fetchQuery_index) begin
        _T_257_218_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_218_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hda == io_fetchQuery_index) begin
        _T_257_218_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_218_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hda == io_fetchQuery_index) begin
        _T_257_218_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_219_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hdb == io_fetchQuery_index) begin
        _T_257_219_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_219_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hdb == io_fetchQuery_index) begin
        _T_257_219_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_219_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hdb == io_fetchQuery_index) begin
        _T_257_219_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_219_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hdb == io_fetchQuery_index) begin
        _T_257_219_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_220_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hdc == io_fetchQuery_index) begin
        _T_257_220_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_220_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hdc == io_fetchQuery_index) begin
        _T_257_220_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_220_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hdc == io_fetchQuery_index) begin
        _T_257_220_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_220_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hdc == io_fetchQuery_index) begin
        _T_257_220_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_221_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hdd == io_fetchQuery_index) begin
        _T_257_221_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_221_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hdd == io_fetchQuery_index) begin
        _T_257_221_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_221_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hdd == io_fetchQuery_index) begin
        _T_257_221_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_221_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hdd == io_fetchQuery_index) begin
        _T_257_221_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_222_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hde == io_fetchQuery_index) begin
        _T_257_222_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_222_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hde == io_fetchQuery_index) begin
        _T_257_222_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_222_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hde == io_fetchQuery_index) begin
        _T_257_222_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_222_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hde == io_fetchQuery_index) begin
        _T_257_222_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_223_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hdf == io_fetchQuery_index) begin
        _T_257_223_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_223_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hdf == io_fetchQuery_index) begin
        _T_257_223_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_223_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hdf == io_fetchQuery_index) begin
        _T_257_223_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_223_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hdf == io_fetchQuery_index) begin
        _T_257_223_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_224_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'he0 == io_fetchQuery_index) begin
        _T_257_224_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_224_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'he0 == io_fetchQuery_index) begin
        _T_257_224_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_224_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'he0 == io_fetchQuery_index) begin
        _T_257_224_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_224_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'he0 == io_fetchQuery_index) begin
        _T_257_224_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_225_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'he1 == io_fetchQuery_index) begin
        _T_257_225_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_225_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'he1 == io_fetchQuery_index) begin
        _T_257_225_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_225_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'he1 == io_fetchQuery_index) begin
        _T_257_225_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_225_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'he1 == io_fetchQuery_index) begin
        _T_257_225_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_226_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'he2 == io_fetchQuery_index) begin
        _T_257_226_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_226_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'he2 == io_fetchQuery_index) begin
        _T_257_226_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_226_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'he2 == io_fetchQuery_index) begin
        _T_257_226_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_226_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'he2 == io_fetchQuery_index) begin
        _T_257_226_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_227_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'he3 == io_fetchQuery_index) begin
        _T_257_227_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_227_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'he3 == io_fetchQuery_index) begin
        _T_257_227_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_227_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'he3 == io_fetchQuery_index) begin
        _T_257_227_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_227_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'he3 == io_fetchQuery_index) begin
        _T_257_227_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_228_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'he4 == io_fetchQuery_index) begin
        _T_257_228_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_228_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'he4 == io_fetchQuery_index) begin
        _T_257_228_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_228_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'he4 == io_fetchQuery_index) begin
        _T_257_228_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_228_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'he4 == io_fetchQuery_index) begin
        _T_257_228_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_229_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'he5 == io_fetchQuery_index) begin
        _T_257_229_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_229_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'he5 == io_fetchQuery_index) begin
        _T_257_229_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_229_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'he5 == io_fetchQuery_index) begin
        _T_257_229_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_229_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'he5 == io_fetchQuery_index) begin
        _T_257_229_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_230_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'he6 == io_fetchQuery_index) begin
        _T_257_230_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_230_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'he6 == io_fetchQuery_index) begin
        _T_257_230_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_230_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'he6 == io_fetchQuery_index) begin
        _T_257_230_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_230_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'he6 == io_fetchQuery_index) begin
        _T_257_230_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_231_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'he7 == io_fetchQuery_index) begin
        _T_257_231_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_231_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'he7 == io_fetchQuery_index) begin
        _T_257_231_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_231_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'he7 == io_fetchQuery_index) begin
        _T_257_231_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_231_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'he7 == io_fetchQuery_index) begin
        _T_257_231_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_232_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'he8 == io_fetchQuery_index) begin
        _T_257_232_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_232_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'he8 == io_fetchQuery_index) begin
        _T_257_232_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_232_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'he8 == io_fetchQuery_index) begin
        _T_257_232_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_232_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'he8 == io_fetchQuery_index) begin
        _T_257_232_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_233_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'he9 == io_fetchQuery_index) begin
        _T_257_233_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_233_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'he9 == io_fetchQuery_index) begin
        _T_257_233_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_233_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'he9 == io_fetchQuery_index) begin
        _T_257_233_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_233_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'he9 == io_fetchQuery_index) begin
        _T_257_233_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_234_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hea == io_fetchQuery_index) begin
        _T_257_234_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_234_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hea == io_fetchQuery_index) begin
        _T_257_234_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_234_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hea == io_fetchQuery_index) begin
        _T_257_234_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_234_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hea == io_fetchQuery_index) begin
        _T_257_234_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_235_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'heb == io_fetchQuery_index) begin
        _T_257_235_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_235_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'heb == io_fetchQuery_index) begin
        _T_257_235_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_235_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'heb == io_fetchQuery_index) begin
        _T_257_235_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_235_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'heb == io_fetchQuery_index) begin
        _T_257_235_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_236_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hec == io_fetchQuery_index) begin
        _T_257_236_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_236_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hec == io_fetchQuery_index) begin
        _T_257_236_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_236_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hec == io_fetchQuery_index) begin
        _T_257_236_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_236_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hec == io_fetchQuery_index) begin
        _T_257_236_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_237_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hed == io_fetchQuery_index) begin
        _T_257_237_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_237_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hed == io_fetchQuery_index) begin
        _T_257_237_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_237_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hed == io_fetchQuery_index) begin
        _T_257_237_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_237_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hed == io_fetchQuery_index) begin
        _T_257_237_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_238_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hee == io_fetchQuery_index) begin
        _T_257_238_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_238_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hee == io_fetchQuery_index) begin
        _T_257_238_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_238_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hee == io_fetchQuery_index) begin
        _T_257_238_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_238_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hee == io_fetchQuery_index) begin
        _T_257_238_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_239_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hef == io_fetchQuery_index) begin
        _T_257_239_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_239_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hef == io_fetchQuery_index) begin
        _T_257_239_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_239_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hef == io_fetchQuery_index) begin
        _T_257_239_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_239_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hef == io_fetchQuery_index) begin
        _T_257_239_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_240_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hf0 == io_fetchQuery_index) begin
        _T_257_240_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_240_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hf0 == io_fetchQuery_index) begin
        _T_257_240_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_240_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hf0 == io_fetchQuery_index) begin
        _T_257_240_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_240_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hf0 == io_fetchQuery_index) begin
        _T_257_240_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_241_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hf1 == io_fetchQuery_index) begin
        _T_257_241_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_241_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hf1 == io_fetchQuery_index) begin
        _T_257_241_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_241_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hf1 == io_fetchQuery_index) begin
        _T_257_241_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_241_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hf1 == io_fetchQuery_index) begin
        _T_257_241_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_242_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hf2 == io_fetchQuery_index) begin
        _T_257_242_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_242_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hf2 == io_fetchQuery_index) begin
        _T_257_242_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_242_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hf2 == io_fetchQuery_index) begin
        _T_257_242_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_242_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hf2 == io_fetchQuery_index) begin
        _T_257_242_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_243_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hf3 == io_fetchQuery_index) begin
        _T_257_243_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_243_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hf3 == io_fetchQuery_index) begin
        _T_257_243_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_243_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hf3 == io_fetchQuery_index) begin
        _T_257_243_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_243_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hf3 == io_fetchQuery_index) begin
        _T_257_243_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_244_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hf4 == io_fetchQuery_index) begin
        _T_257_244_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_244_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hf4 == io_fetchQuery_index) begin
        _T_257_244_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_244_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hf4 == io_fetchQuery_index) begin
        _T_257_244_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_244_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hf4 == io_fetchQuery_index) begin
        _T_257_244_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_245_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hf5 == io_fetchQuery_index) begin
        _T_257_245_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_245_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hf5 == io_fetchQuery_index) begin
        _T_257_245_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_245_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hf5 == io_fetchQuery_index) begin
        _T_257_245_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_245_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hf5 == io_fetchQuery_index) begin
        _T_257_245_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_246_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hf6 == io_fetchQuery_index) begin
        _T_257_246_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_246_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hf6 == io_fetchQuery_index) begin
        _T_257_246_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_246_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hf6 == io_fetchQuery_index) begin
        _T_257_246_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_246_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hf6 == io_fetchQuery_index) begin
        _T_257_246_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_247_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hf7 == io_fetchQuery_index) begin
        _T_257_247_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_247_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hf7 == io_fetchQuery_index) begin
        _T_257_247_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_247_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hf7 == io_fetchQuery_index) begin
        _T_257_247_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_247_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hf7 == io_fetchQuery_index) begin
        _T_257_247_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_248_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hf8 == io_fetchQuery_index) begin
        _T_257_248_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_248_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hf8 == io_fetchQuery_index) begin
        _T_257_248_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_248_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hf8 == io_fetchQuery_index) begin
        _T_257_248_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_248_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hf8 == io_fetchQuery_index) begin
        _T_257_248_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_249_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hf9 == io_fetchQuery_index) begin
        _T_257_249_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_249_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hf9 == io_fetchQuery_index) begin
        _T_257_249_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_249_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hf9 == io_fetchQuery_index) begin
        _T_257_249_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_249_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hf9 == io_fetchQuery_index) begin
        _T_257_249_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_250_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hfa == io_fetchQuery_index) begin
        _T_257_250_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_250_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hfa == io_fetchQuery_index) begin
        _T_257_250_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_250_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hfa == io_fetchQuery_index) begin
        _T_257_250_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_250_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hfa == io_fetchQuery_index) begin
        _T_257_250_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_251_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hfb == io_fetchQuery_index) begin
        _T_257_251_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_251_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hfb == io_fetchQuery_index) begin
        _T_257_251_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_251_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hfb == io_fetchQuery_index) begin
        _T_257_251_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_251_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hfb == io_fetchQuery_index) begin
        _T_257_251_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_252_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hfc == io_fetchQuery_index) begin
        _T_257_252_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_252_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hfc == io_fetchQuery_index) begin
        _T_257_252_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_252_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hfc == io_fetchQuery_index) begin
        _T_257_252_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_252_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hfc == io_fetchQuery_index) begin
        _T_257_252_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_253_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hfd == io_fetchQuery_index) begin
        _T_257_253_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_253_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hfd == io_fetchQuery_index) begin
        _T_257_253_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_253_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hfd == io_fetchQuery_index) begin
        _T_257_253_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_253_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hfd == io_fetchQuery_index) begin
        _T_257_253_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_254_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hfe == io_fetchQuery_index) begin
        _T_257_254_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_254_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hfe == io_fetchQuery_index) begin
        _T_257_254_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_254_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hfe == io_fetchQuery_index) begin
        _T_257_254_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_254_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hfe == io_fetchQuery_index) begin
        _T_257_254_3 <= _T_301_3;
      end
    end
    if (reset) begin
      _T_257_255_0 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hff == io_fetchQuery_index) begin
        _T_257_255_0 <= _T_301_0;
      end
    end
    if (reset) begin
      _T_257_255_1 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hff == io_fetchQuery_index) begin
        _T_257_255_1 <= _T_301_1;
      end
    end
    if (reset) begin
      _T_257_255_2 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hff == io_fetchQuery_index) begin
        _T_257_255_2 <= _T_301_2;
      end
    end
    if (reset) begin
      _T_257_255_3 <= 1'h0;
    end else if (hitInBank) begin
      if (8'hff == io_fetchQuery_index) begin
        _T_257_255_3 <= _T_301_3;
      end
    end
  end
endmodule
module SinglePortBRam(
  input         clock,
  input  [7:0]  io_addr,
  input         io_writeVector,
  input  [31:0] io_inData,
  output [31:0] io_outData
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] _T [0:255]; // @[SinglePortBRam.scala 59:29]
  wire [31:0] _T__T_3_data; // @[SinglePortBRam.scala 59:29]
  wire [7:0] _T__T_3_addr; // @[SinglePortBRam.scala 59:29]
  wire [31:0] _T__T_2_data; // @[SinglePortBRam.scala 59:29]
  wire [7:0] _T__T_2_addr; // @[SinglePortBRam.scala 59:29]
  wire  _T__T_2_mask; // @[SinglePortBRam.scala 59:29]
  wire  _T__T_2_en; // @[SinglePortBRam.scala 59:29]
  reg  _T__T_3_en_pipe_0;
  reg [7:0] _T__T_3_addr_pipe_0;
  assign _T__T_3_addr = _T__T_3_addr_pipe_0;
  assign _T__T_3_data = _T[_T__T_3_addr]; // @[SinglePortBRam.scala 59:29]
  assign _T__T_2_data = io_inData;
  assign _T__T_2_addr = io_addr;
  assign _T__T_2_mask = 1'h1;
  assign _T__T_2_en = io_writeVector;
  assign io_outData = _T__T_3_data; // @[SinglePortBRam.scala 65:22]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    _T[initvar] = _RAND_0[31:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T__T_3_en_pipe_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  _T__T_3_addr_pipe_0 = _RAND_2[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(_T__T_2_en & _T__T_2_mask) begin
      _T[_T__T_2_addr] <= _T__T_2_data; // @[SinglePortBRam.scala 59:29]
    end
    if (io_writeVector) begin
      _T__T_3_en_pipe_0 <= 1'h0;
    end else begin
      _T__T_3_en_pipe_0 <= 1'h1;
    end
    if (io_writeVector ? 1'h0 : 1'h1) begin
      _T__T_3_addr_pipe_0 <= io_addr;
    end
  end
endmodule
module InstBanks(
  input         clock,
  input  [7:0]  io_way_bank_0_0_addr,
  input         io_way_bank_0_0_writeEnable,
  input  [31:0] io_way_bank_0_0_writeData,
  output [31:0] io_way_bank_0_0_readData,
  input  [7:0]  io_way_bank_0_1_addr,
  input         io_way_bank_0_1_writeEnable,
  input  [31:0] io_way_bank_0_1_writeData,
  output [31:0] io_way_bank_0_1_readData,
  input  [7:0]  io_way_bank_1_0_addr,
  input         io_way_bank_1_0_writeEnable,
  input  [31:0] io_way_bank_1_0_writeData,
  output [31:0] io_way_bank_1_0_readData,
  input  [7:0]  io_way_bank_1_1_addr,
  input         io_way_bank_1_1_writeEnable,
  input  [31:0] io_way_bank_1_1_writeData,
  output [31:0] io_way_bank_1_1_readData,
  input  [7:0]  io_way_bank_2_0_addr,
  input         io_way_bank_2_0_writeEnable,
  input  [31:0] io_way_bank_2_0_writeData,
  output [31:0] io_way_bank_2_0_readData,
  input  [7:0]  io_way_bank_2_1_addr,
  input         io_way_bank_2_1_writeEnable,
  input  [31:0] io_way_bank_2_1_writeData,
  output [31:0] io_way_bank_2_1_readData,
  input  [7:0]  io_way_bank_3_0_addr,
  input         io_way_bank_3_0_writeEnable,
  input  [31:0] io_way_bank_3_0_writeData,
  output [31:0] io_way_bank_3_0_readData,
  input  [7:0]  io_way_bank_3_1_addr,
  input         io_way_bank_3_1_writeEnable,
  input  [31:0] io_way_bank_3_1_writeData,
  output [31:0] io_way_bank_3_1_readData
);
  wire  instruction_bank_way_0_bankoffset_0_clock; // @[InstBanks.scala 31:22]
  wire [7:0] instruction_bank_way_0_bankoffset_0_io_addr; // @[InstBanks.scala 31:22]
  wire  instruction_bank_way_0_bankoffset_0_io_writeVector; // @[InstBanks.scala 31:22]
  wire [31:0] instruction_bank_way_0_bankoffset_0_io_inData; // @[InstBanks.scala 31:22]
  wire [31:0] instruction_bank_way_0_bankoffset_0_io_outData; // @[InstBanks.scala 31:22]
  wire  instruction_bank_way_0_bankoffset_1_clock; // @[InstBanks.scala 31:22]
  wire [7:0] instruction_bank_way_0_bankoffset_1_io_addr; // @[InstBanks.scala 31:22]
  wire  instruction_bank_way_0_bankoffset_1_io_writeVector; // @[InstBanks.scala 31:22]
  wire [31:0] instruction_bank_way_0_bankoffset_1_io_inData; // @[InstBanks.scala 31:22]
  wire [31:0] instruction_bank_way_0_bankoffset_1_io_outData; // @[InstBanks.scala 31:22]
  wire  instruction_bank_way_1_bankoffset_0_clock; // @[InstBanks.scala 31:22]
  wire [7:0] instruction_bank_way_1_bankoffset_0_io_addr; // @[InstBanks.scala 31:22]
  wire  instruction_bank_way_1_bankoffset_0_io_writeVector; // @[InstBanks.scala 31:22]
  wire [31:0] instruction_bank_way_1_bankoffset_0_io_inData; // @[InstBanks.scala 31:22]
  wire [31:0] instruction_bank_way_1_bankoffset_0_io_outData; // @[InstBanks.scala 31:22]
  wire  instruction_bank_way_1_bankoffset_1_clock; // @[InstBanks.scala 31:22]
  wire [7:0] instruction_bank_way_1_bankoffset_1_io_addr; // @[InstBanks.scala 31:22]
  wire  instruction_bank_way_1_bankoffset_1_io_writeVector; // @[InstBanks.scala 31:22]
  wire [31:0] instruction_bank_way_1_bankoffset_1_io_inData; // @[InstBanks.scala 31:22]
  wire [31:0] instruction_bank_way_1_bankoffset_1_io_outData; // @[InstBanks.scala 31:22]
  wire  instruction_bank_way_2_bankoffset_0_clock; // @[InstBanks.scala 31:22]
  wire [7:0] instruction_bank_way_2_bankoffset_0_io_addr; // @[InstBanks.scala 31:22]
  wire  instruction_bank_way_2_bankoffset_0_io_writeVector; // @[InstBanks.scala 31:22]
  wire [31:0] instruction_bank_way_2_bankoffset_0_io_inData; // @[InstBanks.scala 31:22]
  wire [31:0] instruction_bank_way_2_bankoffset_0_io_outData; // @[InstBanks.scala 31:22]
  wire  instruction_bank_way_2_bankoffset_1_clock; // @[InstBanks.scala 31:22]
  wire [7:0] instruction_bank_way_2_bankoffset_1_io_addr; // @[InstBanks.scala 31:22]
  wire  instruction_bank_way_2_bankoffset_1_io_writeVector; // @[InstBanks.scala 31:22]
  wire [31:0] instruction_bank_way_2_bankoffset_1_io_inData; // @[InstBanks.scala 31:22]
  wire [31:0] instruction_bank_way_2_bankoffset_1_io_outData; // @[InstBanks.scala 31:22]
  wire  instruction_bank_way_3_bankoffset_0_clock; // @[InstBanks.scala 31:22]
  wire [7:0] instruction_bank_way_3_bankoffset_0_io_addr; // @[InstBanks.scala 31:22]
  wire  instruction_bank_way_3_bankoffset_0_io_writeVector; // @[InstBanks.scala 31:22]
  wire [31:0] instruction_bank_way_3_bankoffset_0_io_inData; // @[InstBanks.scala 31:22]
  wire [31:0] instruction_bank_way_3_bankoffset_0_io_outData; // @[InstBanks.scala 31:22]
  wire  instruction_bank_way_3_bankoffset_1_clock; // @[InstBanks.scala 31:22]
  wire [7:0] instruction_bank_way_3_bankoffset_1_io_addr; // @[InstBanks.scala 31:22]
  wire  instruction_bank_way_3_bankoffset_1_io_writeVector; // @[InstBanks.scala 31:22]
  wire [31:0] instruction_bank_way_3_bankoffset_1_io_inData; // @[InstBanks.scala 31:22]
  wire [31:0] instruction_bank_way_3_bankoffset_1_io_outData; // @[InstBanks.scala 31:22]
  SinglePortBRam instruction_bank_way_0_bankoffset_0 ( // @[InstBanks.scala 31:22]
    .clock(instruction_bank_way_0_bankoffset_0_clock),
    .io_addr(instruction_bank_way_0_bankoffset_0_io_addr),
    .io_writeVector(instruction_bank_way_0_bankoffset_0_io_writeVector),
    .io_inData(instruction_bank_way_0_bankoffset_0_io_inData),
    .io_outData(instruction_bank_way_0_bankoffset_0_io_outData)
  );
  SinglePortBRam instruction_bank_way_0_bankoffset_1 ( // @[InstBanks.scala 31:22]
    .clock(instruction_bank_way_0_bankoffset_1_clock),
    .io_addr(instruction_bank_way_0_bankoffset_1_io_addr),
    .io_writeVector(instruction_bank_way_0_bankoffset_1_io_writeVector),
    .io_inData(instruction_bank_way_0_bankoffset_1_io_inData),
    .io_outData(instruction_bank_way_0_bankoffset_1_io_outData)
  );
  SinglePortBRam instruction_bank_way_1_bankoffset_0 ( // @[InstBanks.scala 31:22]
    .clock(instruction_bank_way_1_bankoffset_0_clock),
    .io_addr(instruction_bank_way_1_bankoffset_0_io_addr),
    .io_writeVector(instruction_bank_way_1_bankoffset_0_io_writeVector),
    .io_inData(instruction_bank_way_1_bankoffset_0_io_inData),
    .io_outData(instruction_bank_way_1_bankoffset_0_io_outData)
  );
  SinglePortBRam instruction_bank_way_1_bankoffset_1 ( // @[InstBanks.scala 31:22]
    .clock(instruction_bank_way_1_bankoffset_1_clock),
    .io_addr(instruction_bank_way_1_bankoffset_1_io_addr),
    .io_writeVector(instruction_bank_way_1_bankoffset_1_io_writeVector),
    .io_inData(instruction_bank_way_1_bankoffset_1_io_inData),
    .io_outData(instruction_bank_way_1_bankoffset_1_io_outData)
  );
  SinglePortBRam instruction_bank_way_2_bankoffset_0 ( // @[InstBanks.scala 31:22]
    .clock(instruction_bank_way_2_bankoffset_0_clock),
    .io_addr(instruction_bank_way_2_bankoffset_0_io_addr),
    .io_writeVector(instruction_bank_way_2_bankoffset_0_io_writeVector),
    .io_inData(instruction_bank_way_2_bankoffset_0_io_inData),
    .io_outData(instruction_bank_way_2_bankoffset_0_io_outData)
  );
  SinglePortBRam instruction_bank_way_2_bankoffset_1 ( // @[InstBanks.scala 31:22]
    .clock(instruction_bank_way_2_bankoffset_1_clock),
    .io_addr(instruction_bank_way_2_bankoffset_1_io_addr),
    .io_writeVector(instruction_bank_way_2_bankoffset_1_io_writeVector),
    .io_inData(instruction_bank_way_2_bankoffset_1_io_inData),
    .io_outData(instruction_bank_way_2_bankoffset_1_io_outData)
  );
  SinglePortBRam instruction_bank_way_3_bankoffset_0 ( // @[InstBanks.scala 31:22]
    .clock(instruction_bank_way_3_bankoffset_0_clock),
    .io_addr(instruction_bank_way_3_bankoffset_0_io_addr),
    .io_writeVector(instruction_bank_way_3_bankoffset_0_io_writeVector),
    .io_inData(instruction_bank_way_3_bankoffset_0_io_inData),
    .io_outData(instruction_bank_way_3_bankoffset_0_io_outData)
  );
  SinglePortBRam instruction_bank_way_3_bankoffset_1 ( // @[InstBanks.scala 31:22]
    .clock(instruction_bank_way_3_bankoffset_1_clock),
    .io_addr(instruction_bank_way_3_bankoffset_1_io_addr),
    .io_writeVector(instruction_bank_way_3_bankoffset_1_io_writeVector),
    .io_inData(instruction_bank_way_3_bankoffset_1_io_inData),
    .io_outData(instruction_bank_way_3_bankoffset_1_io_outData)
  );
  assign io_way_bank_0_0_readData = instruction_bank_way_0_bankoffset_0_io_outData; // @[InstBanks.scala 38:32]
  assign io_way_bank_0_1_readData = instruction_bank_way_0_bankoffset_1_io_outData; // @[InstBanks.scala 38:32]
  assign io_way_bank_1_0_readData = instruction_bank_way_1_bankoffset_0_io_outData; // @[InstBanks.scala 38:32]
  assign io_way_bank_1_1_readData = instruction_bank_way_1_bankoffset_1_io_outData; // @[InstBanks.scala 38:32]
  assign io_way_bank_2_0_readData = instruction_bank_way_2_bankoffset_0_io_outData; // @[InstBanks.scala 38:32]
  assign io_way_bank_2_1_readData = instruction_bank_way_2_bankoffset_1_io_outData; // @[InstBanks.scala 38:32]
  assign io_way_bank_3_0_readData = instruction_bank_way_3_bankoffset_0_io_outData; // @[InstBanks.scala 38:32]
  assign io_way_bank_3_1_readData = instruction_bank_way_3_bankoffset_1_io_outData; // @[InstBanks.scala 38:32]
  assign instruction_bank_way_0_bankoffset_0_clock = clock;
  assign instruction_bank_way_0_bankoffset_0_io_addr = io_way_bank_0_0_addr; // @[InstBanks.scala 35:18]
  assign instruction_bank_way_0_bankoffset_0_io_writeVector = io_way_bank_0_0_writeEnable; // @[InstBanks.scala 37:25]
  assign instruction_bank_way_0_bankoffset_0_io_inData = io_way_bank_0_0_writeData; // @[InstBanks.scala 36:20]
  assign instruction_bank_way_0_bankoffset_1_clock = clock;
  assign instruction_bank_way_0_bankoffset_1_io_addr = io_way_bank_0_1_addr; // @[InstBanks.scala 35:18]
  assign instruction_bank_way_0_bankoffset_1_io_writeVector = io_way_bank_0_1_writeEnable; // @[InstBanks.scala 37:25]
  assign instruction_bank_way_0_bankoffset_1_io_inData = io_way_bank_0_1_writeData; // @[InstBanks.scala 36:20]
  assign instruction_bank_way_1_bankoffset_0_clock = clock;
  assign instruction_bank_way_1_bankoffset_0_io_addr = io_way_bank_1_0_addr; // @[InstBanks.scala 35:18]
  assign instruction_bank_way_1_bankoffset_0_io_writeVector = io_way_bank_1_0_writeEnable; // @[InstBanks.scala 37:25]
  assign instruction_bank_way_1_bankoffset_0_io_inData = io_way_bank_1_0_writeData; // @[InstBanks.scala 36:20]
  assign instruction_bank_way_1_bankoffset_1_clock = clock;
  assign instruction_bank_way_1_bankoffset_1_io_addr = io_way_bank_1_1_addr; // @[InstBanks.scala 35:18]
  assign instruction_bank_way_1_bankoffset_1_io_writeVector = io_way_bank_1_1_writeEnable; // @[InstBanks.scala 37:25]
  assign instruction_bank_way_1_bankoffset_1_io_inData = io_way_bank_1_1_writeData; // @[InstBanks.scala 36:20]
  assign instruction_bank_way_2_bankoffset_0_clock = clock;
  assign instruction_bank_way_2_bankoffset_0_io_addr = io_way_bank_2_0_addr; // @[InstBanks.scala 35:18]
  assign instruction_bank_way_2_bankoffset_0_io_writeVector = io_way_bank_2_0_writeEnable; // @[InstBanks.scala 37:25]
  assign instruction_bank_way_2_bankoffset_0_io_inData = io_way_bank_2_0_writeData; // @[InstBanks.scala 36:20]
  assign instruction_bank_way_2_bankoffset_1_clock = clock;
  assign instruction_bank_way_2_bankoffset_1_io_addr = io_way_bank_2_1_addr; // @[InstBanks.scala 35:18]
  assign instruction_bank_way_2_bankoffset_1_io_writeVector = io_way_bank_2_1_writeEnable; // @[InstBanks.scala 37:25]
  assign instruction_bank_way_2_bankoffset_1_io_inData = io_way_bank_2_1_writeData; // @[InstBanks.scala 36:20]
  assign instruction_bank_way_3_bankoffset_0_clock = clock;
  assign instruction_bank_way_3_bankoffset_0_io_addr = io_way_bank_3_0_addr; // @[InstBanks.scala 35:18]
  assign instruction_bank_way_3_bankoffset_0_io_writeVector = io_way_bank_3_0_writeEnable; // @[InstBanks.scala 37:25]
  assign instruction_bank_way_3_bankoffset_0_io_inData = io_way_bank_3_0_writeData; // @[InstBanks.scala 36:20]
  assign instruction_bank_way_3_bankoffset_1_clock = clock;
  assign instruction_bank_way_3_bankoffset_1_io_addr = io_way_bank_3_1_addr; // @[InstBanks.scala 35:18]
  assign instruction_bank_way_3_bankoffset_1_io_writeVector = io_way_bank_3_1_writeEnable; // @[InstBanks.scala 37:25]
  assign instruction_bank_way_3_bankoffset_1_io_inData = io_way_bank_3_1_writeData; // @[InstBanks.scala 36:20]
endmodule
module ICacheController(
  input   io_flushReq,
  input   io_stage2Free,
  input   io_writeBack,
  output  io_reqReady,
  output  io_writeEnable,
  output  io_flush
);
  wire  _T = ~io_writeBack; // @[ICacheController.scala 36:38]
  assign io_reqReady = io_stage2Free & _T; // @[ICacheController.scala 36:18]
  assign io_writeEnable = io_writeBack; // @[ICacheController.scala 38:18]
  assign io_flush = io_flushReq; // @[ICacheController.scala 37:18]
endmodule
module InstrCache(
  input         clock,
  input         reset,
  output        io_addr_ready,
  input         io_addr_valid,
  input  [31:0] io_addr_bits,
  input         io_data_ready,
  output        io_data_valid,
  output [31:0] io_data_bits,
  input         io_flush,
  input         io_axi_ar_ready,
  output        io_axi_ar_valid,
  output [31:0] io_axi_ar_bits_addr,
  output        io_axi_r_ready,
  input         io_axi_r_valid,
  input  [31:0] io_axi_r_bits_data,
  input         io_axi_r_bits_last
);
  wire  fetch_clock; // @[InstrCache.scala 32:27]
  wire  fetch_reset; // @[InstrCache.scala 32:27]
  wire [31:0] fetch_io_addr; // @[InstrCache.scala 32:27]
  wire  fetch_io_writeTagValid_valid; // @[InstrCache.scala 32:27]
  wire [1:0] fetch_io_writeTagValid_bits_waySelection; // @[InstrCache.scala 32:27]
  wire [7:0] fetch_io_writeTagValid_bits_indexSelection; // @[InstrCache.scala 32:27]
  wire [19:0] fetch_io_writeTagValid_bits_tagValid_tag; // @[InstrCache.scala 32:27]
  wire [7:0] fetch_io_index; // @[InstrCache.scala 32:27]
  wire [19:0] fetch_io_tagValid_0_tag; // @[InstrCache.scala 32:27]
  wire  fetch_io_tagValid_0_valid; // @[InstrCache.scala 32:27]
  wire [19:0] fetch_io_tagValid_1_tag; // @[InstrCache.scala 32:27]
  wire  fetch_io_tagValid_1_valid; // @[InstrCache.scala 32:27]
  wire [19:0] fetch_io_tagValid_2_tag; // @[InstrCache.scala 32:27]
  wire  fetch_io_tagValid_2_valid; // @[InstrCache.scala 32:27]
  wire [19:0] fetch_io_tagValid_3_tag; // @[InstrCache.scala 32:27]
  wire  fetch_io_tagValid_3_valid; // @[InstrCache.scala 32:27]
  wire [19:0] fetch_io_phyTag; // @[InstrCache.scala 32:27]
  wire  fetch_io_bankIndex; // @[InstrCache.scala 32:27]
  wire  fetch_query_clock; // @[InstrCache.scala 33:27]
  wire  fetch_query_reset; // @[InstrCache.scala 33:27]
  wire  fetch_query_io_stall; // @[InstrCache.scala 33:27]
  wire [19:0] fetch_query_io_in_tagValid_0_tag; // @[InstrCache.scala 33:27]
  wire  fetch_query_io_in_tagValid_0_valid; // @[InstrCache.scala 33:27]
  wire [19:0] fetch_query_io_in_tagValid_1_tag; // @[InstrCache.scala 33:27]
  wire  fetch_query_io_in_tagValid_1_valid; // @[InstrCache.scala 33:27]
  wire [19:0] fetch_query_io_in_tagValid_2_tag; // @[InstrCache.scala 33:27]
  wire  fetch_query_io_in_tagValid_2_valid; // @[InstrCache.scala 33:27]
  wire [19:0] fetch_query_io_in_tagValid_3_tag; // @[InstrCache.scala 33:27]
  wire  fetch_query_io_in_tagValid_3_valid; // @[InstrCache.scala 33:27]
  wire [19:0] fetch_query_io_in_phyTag; // @[InstrCache.scala 33:27]
  wire [7:0] fetch_query_io_in_index; // @[InstrCache.scala 33:27]
  wire  fetch_query_io_in_bankIndex; // @[InstrCache.scala 33:27]
  wire  fetch_query_io_in_valid; // @[InstrCache.scala 33:27]
  wire [19:0] fetch_query_io_out_tagValid_0_tag; // @[InstrCache.scala 33:27]
  wire  fetch_query_io_out_tagValid_0_valid; // @[InstrCache.scala 33:27]
  wire [19:0] fetch_query_io_out_tagValid_1_tag; // @[InstrCache.scala 33:27]
  wire  fetch_query_io_out_tagValid_1_valid; // @[InstrCache.scala 33:27]
  wire [19:0] fetch_query_io_out_tagValid_2_tag; // @[InstrCache.scala 33:27]
  wire  fetch_query_io_out_tagValid_2_valid; // @[InstrCache.scala 33:27]
  wire [19:0] fetch_query_io_out_tagValid_3_tag; // @[InstrCache.scala 33:27]
  wire  fetch_query_io_out_tagValid_3_valid; // @[InstrCache.scala 33:27]
  wire [19:0] fetch_query_io_out_phyTag; // @[InstrCache.scala 33:27]
  wire [7:0] fetch_query_io_out_index; // @[InstrCache.scala 33:27]
  wire  fetch_query_io_out_bankIndex; // @[InstrCache.scala 33:27]
  wire  fetch_query_io_out_valid; // @[InstrCache.scala 33:27]
  wire  query_clock; // @[InstrCache.scala 34:27]
  wire  query_reset; // @[InstrCache.scala 34:27]
  wire  query_io_flush; // @[InstrCache.scala 34:27]
  wire  query_io_ready; // @[InstrCache.scala 34:27]
  wire [19:0] query_io_fetchQuery_tagValid_0_tag; // @[InstrCache.scala 34:27]
  wire  query_io_fetchQuery_tagValid_0_valid; // @[InstrCache.scala 34:27]
  wire [19:0] query_io_fetchQuery_tagValid_1_tag; // @[InstrCache.scala 34:27]
  wire  query_io_fetchQuery_tagValid_1_valid; // @[InstrCache.scala 34:27]
  wire [19:0] query_io_fetchQuery_tagValid_2_tag; // @[InstrCache.scala 34:27]
  wire  query_io_fetchQuery_tagValid_2_valid; // @[InstrCache.scala 34:27]
  wire [19:0] query_io_fetchQuery_tagValid_3_tag; // @[InstrCache.scala 34:27]
  wire  query_io_fetchQuery_tagValid_3_valid; // @[InstrCache.scala 34:27]
  wire [19:0] query_io_fetchQuery_phyTag; // @[InstrCache.scala 34:27]
  wire [7:0] query_io_fetchQuery_index; // @[InstrCache.scala 34:27]
  wire  query_io_fetchQuery_bankIndex; // @[InstrCache.scala 34:27]
  wire  query_io_fetchQuery_valid; // @[InstrCache.scala 34:27]
  wire [31:0] query_io_bankData_0; // @[InstrCache.scala 34:27]
  wire [31:0] query_io_bankData_1; // @[InstrCache.scala 34:27]
  wire [31:0] query_io_bankData_2; // @[InstrCache.scala 34:27]
  wire [31:0] query_io_bankData_3; // @[InstrCache.scala 34:27]
  wire  query_io_data_ready; // @[InstrCache.scala 34:27]
  wire  query_io_data_valid; // @[InstrCache.scala 34:27]
  wire [31:0] query_io_data_bits; // @[InstrCache.scala 34:27]
  wire  query_io_writeBundle_writeEnable; // @[InstrCache.scala 34:27]
  wire [1:0] query_io_writeBundle_writeWay; // @[InstrCache.scala 34:27]
  wire [7:0] query_io_writeBundle_writeIndex; // @[InstrCache.scala 34:27]
  wire [19:0] query_io_writeBundle_writeTag; // @[InstrCache.scala 34:27]
  wire [31:0] query_io_writeBundle_writeData_0; // @[InstrCache.scala 34:27]
  wire [31:0] query_io_writeBundle_writeData_1; // @[InstrCache.scala 34:27]
  wire  query_io_axi_ar_ready; // @[InstrCache.scala 34:27]
  wire  query_io_axi_ar_valid; // @[InstrCache.scala 34:27]
  wire [31:0] query_io_axi_ar_bits_addr; // @[InstrCache.scala 34:27]
  wire  query_io_axi_r_ready; // @[InstrCache.scala 34:27]
  wire  query_io_axi_r_valid; // @[InstrCache.scala 34:27]
  wire [31:0] query_io_axi_r_bits_data; // @[InstrCache.scala 34:27]
  wire  query_io_axi_r_bits_last; // @[InstrCache.scala 34:27]
  wire  instrBanks_clock; // @[InstrCache.scala 35:27]
  wire [7:0] instrBanks_io_way_bank_0_0_addr; // @[InstrCache.scala 35:27]
  wire  instrBanks_io_way_bank_0_0_writeEnable; // @[InstrCache.scala 35:27]
  wire [31:0] instrBanks_io_way_bank_0_0_writeData; // @[InstrCache.scala 35:27]
  wire [31:0] instrBanks_io_way_bank_0_0_readData; // @[InstrCache.scala 35:27]
  wire [7:0] instrBanks_io_way_bank_0_1_addr; // @[InstrCache.scala 35:27]
  wire  instrBanks_io_way_bank_0_1_writeEnable; // @[InstrCache.scala 35:27]
  wire [31:0] instrBanks_io_way_bank_0_1_writeData; // @[InstrCache.scala 35:27]
  wire [31:0] instrBanks_io_way_bank_0_1_readData; // @[InstrCache.scala 35:27]
  wire [7:0] instrBanks_io_way_bank_1_0_addr; // @[InstrCache.scala 35:27]
  wire  instrBanks_io_way_bank_1_0_writeEnable; // @[InstrCache.scala 35:27]
  wire [31:0] instrBanks_io_way_bank_1_0_writeData; // @[InstrCache.scala 35:27]
  wire [31:0] instrBanks_io_way_bank_1_0_readData; // @[InstrCache.scala 35:27]
  wire [7:0] instrBanks_io_way_bank_1_1_addr; // @[InstrCache.scala 35:27]
  wire  instrBanks_io_way_bank_1_1_writeEnable; // @[InstrCache.scala 35:27]
  wire [31:0] instrBanks_io_way_bank_1_1_writeData; // @[InstrCache.scala 35:27]
  wire [31:0] instrBanks_io_way_bank_1_1_readData; // @[InstrCache.scala 35:27]
  wire [7:0] instrBanks_io_way_bank_2_0_addr; // @[InstrCache.scala 35:27]
  wire  instrBanks_io_way_bank_2_0_writeEnable; // @[InstrCache.scala 35:27]
  wire [31:0] instrBanks_io_way_bank_2_0_writeData; // @[InstrCache.scala 35:27]
  wire [31:0] instrBanks_io_way_bank_2_0_readData; // @[InstrCache.scala 35:27]
  wire [7:0] instrBanks_io_way_bank_2_1_addr; // @[InstrCache.scala 35:27]
  wire  instrBanks_io_way_bank_2_1_writeEnable; // @[InstrCache.scala 35:27]
  wire [31:0] instrBanks_io_way_bank_2_1_writeData; // @[InstrCache.scala 35:27]
  wire [31:0] instrBanks_io_way_bank_2_1_readData; // @[InstrCache.scala 35:27]
  wire [7:0] instrBanks_io_way_bank_3_0_addr; // @[InstrCache.scala 35:27]
  wire  instrBanks_io_way_bank_3_0_writeEnable; // @[InstrCache.scala 35:27]
  wire [31:0] instrBanks_io_way_bank_3_0_writeData; // @[InstrCache.scala 35:27]
  wire [31:0] instrBanks_io_way_bank_3_0_readData; // @[InstrCache.scala 35:27]
  wire [7:0] instrBanks_io_way_bank_3_1_addr; // @[InstrCache.scala 35:27]
  wire  instrBanks_io_way_bank_3_1_writeEnable; // @[InstrCache.scala 35:27]
  wire [31:0] instrBanks_io_way_bank_3_1_writeData; // @[InstrCache.scala 35:27]
  wire [31:0] instrBanks_io_way_bank_3_1_readData; // @[InstrCache.scala 35:27]
  wire  controller_io_flushReq; // @[InstrCache.scala 36:27]
  wire  controller_io_stage2Free; // @[InstrCache.scala 36:27]
  wire  controller_io_writeBack; // @[InstrCache.scala 36:27]
  wire  controller_io_reqReady; // @[InstrCache.scala 36:27]
  wire  controller_io_writeEnable; // @[InstrCache.scala 36:27]
  wire  controller_io_flush; // @[InstrCache.scala 36:27]
  wire  _T_11 = 2'h0 == query_io_writeBundle_writeWay; // @[InstrCache.scala 63:42]
  wire [31:0] _GEN_3 = instrBanks_io_way_bank_0_0_readData; // @[InstrCache.scala 66:23]
  wire  _T_17 = 2'h1 == query_io_writeBundle_writeWay; // @[InstrCache.scala 63:42]
  wire [31:0] _GEN_11 = instrBanks_io_way_bank_1_0_readData; // @[InstrCache.scala 66:23]
  wire  _T_23 = 2'h2 == query_io_writeBundle_writeWay; // @[InstrCache.scala 63:42]
  wire [31:0] _GEN_19 = instrBanks_io_way_bank_2_0_readData; // @[InstrCache.scala 66:23]
  wire  _T_29 = 2'h3 == query_io_writeBundle_writeWay; // @[InstrCache.scala 63:42]
  wire [31:0] _GEN_27 = instrBanks_io_way_bank_3_0_readData; // @[InstrCache.scala 66:23]
  FetchTop fetch ( // @[InstrCache.scala 32:27]
    .clock(fetch_clock),
    .reset(fetch_reset),
    .io_addr(fetch_io_addr),
    .io_writeTagValid_valid(fetch_io_writeTagValid_valid),
    .io_writeTagValid_bits_waySelection(fetch_io_writeTagValid_bits_waySelection),
    .io_writeTagValid_bits_indexSelection(fetch_io_writeTagValid_bits_indexSelection),
    .io_writeTagValid_bits_tagValid_tag(fetch_io_writeTagValid_bits_tagValid_tag),
    .io_index(fetch_io_index),
    .io_tagValid_0_tag(fetch_io_tagValid_0_tag),
    .io_tagValid_0_valid(fetch_io_tagValid_0_valid),
    .io_tagValid_1_tag(fetch_io_tagValid_1_tag),
    .io_tagValid_1_valid(fetch_io_tagValid_1_valid),
    .io_tagValid_2_tag(fetch_io_tagValid_2_tag),
    .io_tagValid_2_valid(fetch_io_tagValid_2_valid),
    .io_tagValid_3_tag(fetch_io_tagValid_3_tag),
    .io_tagValid_3_valid(fetch_io_tagValid_3_valid),
    .io_phyTag(fetch_io_phyTag),
    .io_bankIndex(fetch_io_bankIndex)
  );
  CachePipelineStage fetch_query ( // @[InstrCache.scala 33:27]
    .clock(fetch_query_clock),
    .reset(fetch_query_reset),
    .io_stall(fetch_query_io_stall),
    .io_in_tagValid_0_tag(fetch_query_io_in_tagValid_0_tag),
    .io_in_tagValid_0_valid(fetch_query_io_in_tagValid_0_valid),
    .io_in_tagValid_1_tag(fetch_query_io_in_tagValid_1_tag),
    .io_in_tagValid_1_valid(fetch_query_io_in_tagValid_1_valid),
    .io_in_tagValid_2_tag(fetch_query_io_in_tagValid_2_tag),
    .io_in_tagValid_2_valid(fetch_query_io_in_tagValid_2_valid),
    .io_in_tagValid_3_tag(fetch_query_io_in_tagValid_3_tag),
    .io_in_tagValid_3_valid(fetch_query_io_in_tagValid_3_valid),
    .io_in_phyTag(fetch_query_io_in_phyTag),
    .io_in_index(fetch_query_io_in_index),
    .io_in_bankIndex(fetch_query_io_in_bankIndex),
    .io_in_valid(fetch_query_io_in_valid),
    .io_out_tagValid_0_tag(fetch_query_io_out_tagValid_0_tag),
    .io_out_tagValid_0_valid(fetch_query_io_out_tagValid_0_valid),
    .io_out_tagValid_1_tag(fetch_query_io_out_tagValid_1_tag),
    .io_out_tagValid_1_valid(fetch_query_io_out_tagValid_1_valid),
    .io_out_tagValid_2_tag(fetch_query_io_out_tagValid_2_tag),
    .io_out_tagValid_2_valid(fetch_query_io_out_tagValid_2_valid),
    .io_out_tagValid_3_tag(fetch_query_io_out_tagValid_3_tag),
    .io_out_tagValid_3_valid(fetch_query_io_out_tagValid_3_valid),
    .io_out_phyTag(fetch_query_io_out_phyTag),
    .io_out_index(fetch_query_io_out_index),
    .io_out_bankIndex(fetch_query_io_out_bankIndex),
    .io_out_valid(fetch_query_io_out_valid)
  );
  QueryTop query ( // @[InstrCache.scala 34:27]
    .clock(query_clock),
    .reset(query_reset),
    .io_flush(query_io_flush),
    .io_ready(query_io_ready),
    .io_fetchQuery_tagValid_0_tag(query_io_fetchQuery_tagValid_0_tag),
    .io_fetchQuery_tagValid_0_valid(query_io_fetchQuery_tagValid_0_valid),
    .io_fetchQuery_tagValid_1_tag(query_io_fetchQuery_tagValid_1_tag),
    .io_fetchQuery_tagValid_1_valid(query_io_fetchQuery_tagValid_1_valid),
    .io_fetchQuery_tagValid_2_tag(query_io_fetchQuery_tagValid_2_tag),
    .io_fetchQuery_tagValid_2_valid(query_io_fetchQuery_tagValid_2_valid),
    .io_fetchQuery_tagValid_3_tag(query_io_fetchQuery_tagValid_3_tag),
    .io_fetchQuery_tagValid_3_valid(query_io_fetchQuery_tagValid_3_valid),
    .io_fetchQuery_phyTag(query_io_fetchQuery_phyTag),
    .io_fetchQuery_index(query_io_fetchQuery_index),
    .io_fetchQuery_bankIndex(query_io_fetchQuery_bankIndex),
    .io_fetchQuery_valid(query_io_fetchQuery_valid),
    .io_bankData_0(query_io_bankData_0),
    .io_bankData_1(query_io_bankData_1),
    .io_bankData_2(query_io_bankData_2),
    .io_bankData_3(query_io_bankData_3),
    .io_data_ready(query_io_data_ready),
    .io_data_valid(query_io_data_valid),
    .io_data_bits(query_io_data_bits),
    .io_writeBundle_writeEnable(query_io_writeBundle_writeEnable),
    .io_writeBundle_writeWay(query_io_writeBundle_writeWay),
    .io_writeBundle_writeIndex(query_io_writeBundle_writeIndex),
    .io_writeBundle_writeTag(query_io_writeBundle_writeTag),
    .io_writeBundle_writeData_0(query_io_writeBundle_writeData_0),
    .io_writeBundle_writeData_1(query_io_writeBundle_writeData_1),
    .io_axi_ar_ready(query_io_axi_ar_ready),
    .io_axi_ar_valid(query_io_axi_ar_valid),
    .io_axi_ar_bits_addr(query_io_axi_ar_bits_addr),
    .io_axi_r_ready(query_io_axi_r_ready),
    .io_axi_r_valid(query_io_axi_r_valid),
    .io_axi_r_bits_data(query_io_axi_r_bits_data),
    .io_axi_r_bits_last(query_io_axi_r_bits_last)
  );
  InstBanks instrBanks ( // @[InstrCache.scala 35:27]
    .clock(instrBanks_clock),
    .io_way_bank_0_0_addr(instrBanks_io_way_bank_0_0_addr),
    .io_way_bank_0_0_writeEnable(instrBanks_io_way_bank_0_0_writeEnable),
    .io_way_bank_0_0_writeData(instrBanks_io_way_bank_0_0_writeData),
    .io_way_bank_0_0_readData(instrBanks_io_way_bank_0_0_readData),
    .io_way_bank_0_1_addr(instrBanks_io_way_bank_0_1_addr),
    .io_way_bank_0_1_writeEnable(instrBanks_io_way_bank_0_1_writeEnable),
    .io_way_bank_0_1_writeData(instrBanks_io_way_bank_0_1_writeData),
    .io_way_bank_0_1_readData(instrBanks_io_way_bank_0_1_readData),
    .io_way_bank_1_0_addr(instrBanks_io_way_bank_1_0_addr),
    .io_way_bank_1_0_writeEnable(instrBanks_io_way_bank_1_0_writeEnable),
    .io_way_bank_1_0_writeData(instrBanks_io_way_bank_1_0_writeData),
    .io_way_bank_1_0_readData(instrBanks_io_way_bank_1_0_readData),
    .io_way_bank_1_1_addr(instrBanks_io_way_bank_1_1_addr),
    .io_way_bank_1_1_writeEnable(instrBanks_io_way_bank_1_1_writeEnable),
    .io_way_bank_1_1_writeData(instrBanks_io_way_bank_1_1_writeData),
    .io_way_bank_1_1_readData(instrBanks_io_way_bank_1_1_readData),
    .io_way_bank_2_0_addr(instrBanks_io_way_bank_2_0_addr),
    .io_way_bank_2_0_writeEnable(instrBanks_io_way_bank_2_0_writeEnable),
    .io_way_bank_2_0_writeData(instrBanks_io_way_bank_2_0_writeData),
    .io_way_bank_2_0_readData(instrBanks_io_way_bank_2_0_readData),
    .io_way_bank_2_1_addr(instrBanks_io_way_bank_2_1_addr),
    .io_way_bank_2_1_writeEnable(instrBanks_io_way_bank_2_1_writeEnable),
    .io_way_bank_2_1_writeData(instrBanks_io_way_bank_2_1_writeData),
    .io_way_bank_2_1_readData(instrBanks_io_way_bank_2_1_readData),
    .io_way_bank_3_0_addr(instrBanks_io_way_bank_3_0_addr),
    .io_way_bank_3_0_writeEnable(instrBanks_io_way_bank_3_0_writeEnable),
    .io_way_bank_3_0_writeData(instrBanks_io_way_bank_3_0_writeData),
    .io_way_bank_3_0_readData(instrBanks_io_way_bank_3_0_readData),
    .io_way_bank_3_1_addr(instrBanks_io_way_bank_3_1_addr),
    .io_way_bank_3_1_writeEnable(instrBanks_io_way_bank_3_1_writeEnable),
    .io_way_bank_3_1_writeData(instrBanks_io_way_bank_3_1_writeData),
    .io_way_bank_3_1_readData(instrBanks_io_way_bank_3_1_readData)
  );
  ICacheController controller ( // @[InstrCache.scala 36:27]
    .io_flushReq(controller_io_flushReq),
    .io_stage2Free(controller_io_stage2Free),
    .io_writeBack(controller_io_writeBack),
    .io_reqReady(controller_io_reqReady),
    .io_writeEnable(controller_io_writeEnable),
    .io_flush(controller_io_flush)
  );
  assign io_addr_ready = controller_io_reqReady; // @[InstrCache.scala 38:28]
  assign io_data_valid = query_io_data_valid; // @[InstrCache.scala 87:23]
  assign io_data_bits = query_io_data_bits; // @[InstrCache.scala 87:23]
  assign io_axi_ar_valid = query_io_axi_ar_valid; // @[InstrCache.scala 88:23]
  assign io_axi_ar_bits_addr = query_io_axi_ar_bits_addr; // @[InstrCache.scala 88:23]
  assign io_axi_r_ready = query_io_axi_r_ready; // @[InstrCache.scala 88:23]
  assign fetch_clock = clock;
  assign fetch_reset = reset;
  assign fetch_io_addr = io_addr_bits; // @[InstrCache.scala 41:46]
  assign fetch_io_writeTagValid_valid = controller_io_writeEnable; // @[InstrCache.scala 42:46]
  assign fetch_io_writeTagValid_bits_waySelection = query_io_writeBundle_writeWay; // @[InstrCache.scala 50:44]
  assign fetch_io_writeTagValid_bits_indexSelection = query_io_writeBundle_writeIndex; // @[InstrCache.scala 45:46]
  assign fetch_io_writeTagValid_bits_tagValid_tag = query_io_writeBundle_writeTag; // @[InstrCache.scala 43:46]
  assign fetch_query_clock = clock;
  assign fetch_query_reset = reset;
  assign fetch_query_io_stall = ~controller_io_stage2Free; // @[InstrCache.scala 73:31]
  assign fetch_query_io_in_tagValid_0_tag = fetch_io_tagValid_0_tag; // @[InstrCache.scala 75:31]
  assign fetch_query_io_in_tagValid_0_valid = fetch_io_tagValid_0_valid; // @[InstrCache.scala 75:31]
  assign fetch_query_io_in_tagValid_1_tag = fetch_io_tagValid_1_tag; // @[InstrCache.scala 75:31]
  assign fetch_query_io_in_tagValid_1_valid = fetch_io_tagValid_1_valid; // @[InstrCache.scala 75:31]
  assign fetch_query_io_in_tagValid_2_tag = fetch_io_tagValid_2_tag; // @[InstrCache.scala 75:31]
  assign fetch_query_io_in_tagValid_2_valid = fetch_io_tagValid_2_valid; // @[InstrCache.scala 75:31]
  assign fetch_query_io_in_tagValid_3_tag = fetch_io_tagValid_3_tag; // @[InstrCache.scala 75:31]
  assign fetch_query_io_in_tagValid_3_valid = fetch_io_tagValid_3_valid; // @[InstrCache.scala 75:31]
  assign fetch_query_io_in_phyTag = fetch_io_phyTag; // @[InstrCache.scala 76:31]
  assign fetch_query_io_in_index = fetch_io_index; // @[InstrCache.scala 74:31]
  assign fetch_query_io_in_bankIndex = fetch_io_bankIndex; // @[InstrCache.scala 77:31]
  assign fetch_query_io_in_valid = io_addr_ready & io_addr_valid; // @[InstrCache.scala 78:31]
  assign query_clock = clock;
  assign query_reset = reset;
  assign query_io_flush = controller_io_flush; // @[InstrCache.scala 84:23]
  assign query_io_fetchQuery_tagValid_0_tag = fetch_query_io_out_tagValid_0_tag; // @[InstrCache.scala 85:23]
  assign query_io_fetchQuery_tagValid_0_valid = fetch_query_io_out_tagValid_0_valid; // @[InstrCache.scala 85:23]
  assign query_io_fetchQuery_tagValid_1_tag = fetch_query_io_out_tagValid_1_tag; // @[InstrCache.scala 85:23]
  assign query_io_fetchQuery_tagValid_1_valid = fetch_query_io_out_tagValid_1_valid; // @[InstrCache.scala 85:23]
  assign query_io_fetchQuery_tagValid_2_tag = fetch_query_io_out_tagValid_2_tag; // @[InstrCache.scala 85:23]
  assign query_io_fetchQuery_tagValid_2_valid = fetch_query_io_out_tagValid_2_valid; // @[InstrCache.scala 85:23]
  assign query_io_fetchQuery_tagValid_3_tag = fetch_query_io_out_tagValid_3_tag; // @[InstrCache.scala 85:23]
  assign query_io_fetchQuery_tagValid_3_valid = fetch_query_io_out_tagValid_3_valid; // @[InstrCache.scala 85:23]
  assign query_io_fetchQuery_phyTag = fetch_query_io_out_phyTag; // @[InstrCache.scala 85:23]
  assign query_io_fetchQuery_index = fetch_query_io_out_index; // @[InstrCache.scala 85:23]
  assign query_io_fetchQuery_bankIndex = fetch_query_io_out_bankIndex; // @[InstrCache.scala 85:23]
  assign query_io_fetchQuery_valid = fetch_query_io_out_valid; // @[InstrCache.scala 85:23]
  assign query_io_bankData_0 = fetch_query_io_out_bankIndex ? instrBanks_io_way_bank_0_1_readData : _GEN_3; // @[InstrCache.scala 86:23]
  assign query_io_bankData_1 = fetch_query_io_out_bankIndex ? instrBanks_io_way_bank_1_1_readData : _GEN_11; // @[InstrCache.scala 86:23]
  assign query_io_bankData_2 = fetch_query_io_out_bankIndex ? instrBanks_io_way_bank_2_1_readData : _GEN_19; // @[InstrCache.scala 86:23]
  assign query_io_bankData_3 = fetch_query_io_out_bankIndex ? instrBanks_io_way_bank_3_1_readData : _GEN_27; // @[InstrCache.scala 86:23]
  assign query_io_data_ready = io_data_ready; // @[InstrCache.scala 87:23]
  assign query_io_axi_ar_ready = io_axi_ar_ready; // @[InstrCache.scala 88:23]
  assign query_io_axi_r_valid = io_axi_r_valid; // @[InstrCache.scala 88:23]
  assign query_io_axi_r_bits_data = io_axi_r_bits_data; // @[InstrCache.scala 88:23]
  assign query_io_axi_r_bits_last = io_axi_r_bits_last; // @[InstrCache.scala 88:23]
  assign instrBanks_clock = clock;
  assign instrBanks_io_way_bank_0_0_addr = controller_io_writeEnable ? query_io_writeBundle_writeIndex : fetch_io_index; // @[InstrCache.scala 57:41]
  assign instrBanks_io_way_bank_0_0_writeEnable = controller_io_writeEnable & _T_11; // @[InstrCache.scala 62:48]
  assign instrBanks_io_way_bank_0_0_writeData = query_io_writeBundle_writeData_0; // @[InstrCache.scala 64:46]
  assign instrBanks_io_way_bank_0_1_addr = controller_io_writeEnable ? query_io_writeBundle_writeIndex : fetch_io_index; // @[InstrCache.scala 57:41]
  assign instrBanks_io_way_bank_0_1_writeEnable = controller_io_writeEnable & _T_11; // @[InstrCache.scala 62:48]
  assign instrBanks_io_way_bank_0_1_writeData = query_io_writeBundle_writeData_1; // @[InstrCache.scala 64:46]
  assign instrBanks_io_way_bank_1_0_addr = controller_io_writeEnable ? query_io_writeBundle_writeIndex : fetch_io_index; // @[InstrCache.scala 57:41]
  assign instrBanks_io_way_bank_1_0_writeEnable = controller_io_writeEnable & _T_17; // @[InstrCache.scala 62:48]
  assign instrBanks_io_way_bank_1_0_writeData = query_io_writeBundle_writeData_0; // @[InstrCache.scala 64:46]
  assign instrBanks_io_way_bank_1_1_addr = controller_io_writeEnable ? query_io_writeBundle_writeIndex : fetch_io_index; // @[InstrCache.scala 57:41]
  assign instrBanks_io_way_bank_1_1_writeEnable = controller_io_writeEnable & _T_17; // @[InstrCache.scala 62:48]
  assign instrBanks_io_way_bank_1_1_writeData = query_io_writeBundle_writeData_1; // @[InstrCache.scala 64:46]
  assign instrBanks_io_way_bank_2_0_addr = controller_io_writeEnable ? query_io_writeBundle_writeIndex : fetch_io_index; // @[InstrCache.scala 57:41]
  assign instrBanks_io_way_bank_2_0_writeEnable = controller_io_writeEnable & _T_23; // @[InstrCache.scala 62:48]
  assign instrBanks_io_way_bank_2_0_writeData = query_io_writeBundle_writeData_0; // @[InstrCache.scala 64:46]
  assign instrBanks_io_way_bank_2_1_addr = controller_io_writeEnable ? query_io_writeBundle_writeIndex : fetch_io_index; // @[InstrCache.scala 57:41]
  assign instrBanks_io_way_bank_2_1_writeEnable = controller_io_writeEnable & _T_23; // @[InstrCache.scala 62:48]
  assign instrBanks_io_way_bank_2_1_writeData = query_io_writeBundle_writeData_1; // @[InstrCache.scala 64:46]
  assign instrBanks_io_way_bank_3_0_addr = controller_io_writeEnable ? query_io_writeBundle_writeIndex : fetch_io_index; // @[InstrCache.scala 57:41]
  assign instrBanks_io_way_bank_3_0_writeEnable = controller_io_writeEnable & _T_29; // @[InstrCache.scala 62:48]
  assign instrBanks_io_way_bank_3_0_writeData = query_io_writeBundle_writeData_0; // @[InstrCache.scala 64:46]
  assign instrBanks_io_way_bank_3_1_addr = controller_io_writeEnable ? query_io_writeBundle_writeIndex : fetch_io_index; // @[InstrCache.scala 57:41]
  assign instrBanks_io_way_bank_3_1_writeEnable = controller_io_writeEnable & _T_29; // @[InstrCache.scala 62:48]
  assign instrBanks_io_way_bank_3_1_writeData = query_io_writeBundle_writeData_1; // @[InstrCache.scala 64:46]
  assign controller_io_flushReq = io_flush; // @[InstrCache.scala 90:28]
  assign controller_io_stage2Free = query_io_ready; // @[InstrCache.scala 91:28]
  assign controller_io_writeBack = query_io_writeBundle_writeEnable; // @[InstrCache.scala 92:28]
endmodule
module Queue(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [31:0] io_enq_bits_addr,
  input  [3:0]  io_enq_bits_len,
  input  [1:0]  io_enq_bits_burst,
  input         io_deq_ready,
  output        io_deq_valid,
  output [31:0] io_deq_bits_addr,
  output [3:0]  io_deq_bits_len,
  output [1:0]  io_deq_bits_burst
);
`ifdef RANDOMIZE_GARBAGE_ASSIGN
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_5;
`endif // RANDOMIZE_GARBAGE_ASSIGN
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] ram_addr [0:9]; // @[Decoupled.scala 209:16]
  wire [31:0] ram_addr__T_15_data; // @[Decoupled.scala 209:16]
  wire [3:0] ram_addr__T_15_addr; // @[Decoupled.scala 209:16]
  wire [31:0] ram_addr__T_5_data; // @[Decoupled.scala 209:16]
  wire [3:0] ram_addr__T_5_addr; // @[Decoupled.scala 209:16]
  wire  ram_addr__T_5_mask; // @[Decoupled.scala 209:16]
  wire  ram_addr__T_5_en; // @[Decoupled.scala 209:16]
  reg [3:0] ram_len [0:9]; // @[Decoupled.scala 209:16]
  wire [3:0] ram_len__T_15_data; // @[Decoupled.scala 209:16]
  wire [3:0] ram_len__T_15_addr; // @[Decoupled.scala 209:16]
  wire [3:0] ram_len__T_5_data; // @[Decoupled.scala 209:16]
  wire [3:0] ram_len__T_5_addr; // @[Decoupled.scala 209:16]
  wire  ram_len__T_5_mask; // @[Decoupled.scala 209:16]
  wire  ram_len__T_5_en; // @[Decoupled.scala 209:16]
  reg [1:0] ram_burst [0:9]; // @[Decoupled.scala 209:16]
  wire [1:0] ram_burst__T_15_data; // @[Decoupled.scala 209:16]
  wire [3:0] ram_burst__T_15_addr; // @[Decoupled.scala 209:16]
  wire [1:0] ram_burst__T_5_data; // @[Decoupled.scala 209:16]
  wire [3:0] ram_burst__T_5_addr; // @[Decoupled.scala 209:16]
  wire  ram_burst__T_5_mask; // @[Decoupled.scala 209:16]
  wire  ram_burst__T_5_en; // @[Decoupled.scala 209:16]
  reg [3:0] _T; // @[Counter.scala 29:33]
  reg [3:0] _T_1; // @[Counter.scala 29:33]
  reg  maybe_full; // @[Decoupled.scala 212:27]
  wire  ptr_match = _T == _T_1; // @[Decoupled.scala 214:33]
  wire  _T_2 = ~maybe_full; // @[Decoupled.scala 215:28]
  wire  empty = ptr_match & _T_2; // @[Decoupled.scala 215:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 216:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  wire  _T_6 = _T == 4'h9; // @[Counter.scala 38:24]
  wire [3:0] _T_8 = _T + 4'h1; // @[Counter.scala 39:22]
  wire  _T_9 = _T_1 == 4'h9; // @[Counter.scala 38:24]
  wire [3:0] _T_11 = _T_1 + 4'h1; // @[Counter.scala 39:22]
  wire  _T_12 = do_enq != do_deq; // @[Decoupled.scala 227:16]
  assign ram_addr__T_15_addr = _T_1;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_addr__T_15_data = ram_addr[ram_addr__T_15_addr]; // @[Decoupled.scala 209:16]
  `else
  assign ram_addr__T_15_data = ram_addr__T_15_addr >= 4'ha ? _RAND_1[31:0] : ram_addr[ram_addr__T_15_addr]; // @[Decoupled.scala 209:16]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_addr__T_5_data = io_enq_bits_addr;
  assign ram_addr__T_5_addr = _T;
  assign ram_addr__T_5_mask = 1'h1;
  assign ram_addr__T_5_en = io_enq_ready & io_enq_valid;
  assign ram_len__T_15_addr = _T_1;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_len__T_15_data = ram_len[ram_len__T_15_addr]; // @[Decoupled.scala 209:16]
  `else
  assign ram_len__T_15_data = ram_len__T_15_addr >= 4'ha ? _RAND_3[3:0] : ram_len[ram_len__T_15_addr]; // @[Decoupled.scala 209:16]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_len__T_5_data = io_enq_bits_len;
  assign ram_len__T_5_addr = _T;
  assign ram_len__T_5_mask = 1'h1;
  assign ram_len__T_5_en = io_enq_ready & io_enq_valid;
  assign ram_burst__T_15_addr = _T_1;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_burst__T_15_data = ram_burst[ram_burst__T_15_addr]; // @[Decoupled.scala 209:16]
  `else
  assign ram_burst__T_15_data = ram_burst__T_15_addr >= 4'ha ? _RAND_5[1:0] : ram_burst[ram_burst__T_15_addr]; // @[Decoupled.scala 209:16]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_burst__T_5_data = io_enq_bits_burst;
  assign ram_burst__T_5_addr = _T;
  assign ram_burst__T_5_mask = 1'h1;
  assign ram_burst__T_5_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 232:16]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 231:16]
  assign io_deq_bits_addr = ram_addr__T_15_data; // @[Decoupled.scala 233:15]
  assign io_deq_bits_len = ram_len__T_15_data; // @[Decoupled.scala 233:15]
  assign io_deq_bits_burst = ram_burst__T_15_data; // @[Decoupled.scala 233:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_GARBAGE_ASSIGN
  _RAND_1 = {1{`RANDOM}};
  _RAND_3 = {1{`RANDOM}};
  _RAND_5 = {1{`RANDOM}};
`endif // RANDOMIZE_GARBAGE_ASSIGN
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 10; initvar = initvar+1)
    ram_addr[initvar] = _RAND_0[31:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 10; initvar = initvar+1)
    ram_len[initvar] = _RAND_2[3:0];
  _RAND_4 = {1{`RANDOM}};
  for (initvar = 0; initvar < 10; initvar = initvar+1)
    ram_burst[initvar] = _RAND_4[1:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T = _RAND_6[3:0];
  _RAND_7 = {1{`RANDOM}};
  _T_1 = _RAND_7[3:0];
  _RAND_8 = {1{`RANDOM}};
  maybe_full = _RAND_8[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(ram_addr__T_5_en & ram_addr__T_5_mask) begin
      ram_addr[ram_addr__T_5_addr] <= ram_addr__T_5_data; // @[Decoupled.scala 209:16]
    end
    if(ram_len__T_5_en & ram_len__T_5_mask) begin
      ram_len[ram_len__T_5_addr] <= ram_len__T_5_data; // @[Decoupled.scala 209:16]
    end
    if(ram_burst__T_5_en & ram_burst__T_5_mask) begin
      ram_burst[ram_burst__T_5_addr] <= ram_burst__T_5_data; // @[Decoupled.scala 209:16]
    end
    if (reset) begin
      _T <= 4'h0;
    end else if (do_enq) begin
      if (_T_6) begin
        _T <= 4'h0;
      end else begin
        _T <= _T_8;
      end
    end
    if (reset) begin
      _T_1 <= 4'h0;
    end else if (do_deq) begin
      if (_T_9) begin
        _T_1 <= 4'h0;
      end else begin
        _T_1 <= _T_11;
      end
    end
    if (reset) begin
      maybe_full <= 1'h0;
    end else if (_T_12) begin
      maybe_full <= do_enq;
    end
  end
endmodule
module VeriAXIRam(
  input         clock,
  input         reset,
  output        io_axi_ar_ready,
  input         io_axi_ar_valid,
  input  [31:0] io_axi_ar_bits_addr,
  input         io_axi_r_ready,
  output        io_axi_r_valid,
  output [31:0] io_axi_r_bits_data,
  output        io_axi_r_bits_last
);
`ifdef RANDOMIZE_GARBAGE_ASSIGN
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_GARBAGE_ASSIGN
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] mem [0:4094]; // @[VeriAXIRam.scala 21:16]
  wire [31:0] mem__T_92_data; // @[VeriAXIRam.scala 21:16]
  wire [11:0] mem__T_92_addr; // @[VeriAXIRam.scala 21:16]
  wire [31:0] mem_internalData_data; // @[VeriAXIRam.scala 21:16]
  wire [11:0] mem_internalData_addr; // @[VeriAXIRam.scala 21:16]
  wire [31:0] mem__T_155_data; // @[VeriAXIRam.scala 21:16]
  wire [11:0] mem__T_155_addr; // @[VeriAXIRam.scala 21:16]
  wire  mem__T_155_mask; // @[VeriAXIRam.scala 21:16]
  wire  mem__T_155_en; // @[VeriAXIRam.scala 21:16]
  wire  instRQ_clock; // @[VeriAXIRam.scala 34:22]
  wire  instRQ_reset; // @[VeriAXIRam.scala 34:22]
  wire  instRQ_io_enq_ready; // @[VeriAXIRam.scala 34:22]
  wire  instRQ_io_enq_valid; // @[VeriAXIRam.scala 34:22]
  wire [31:0] instRQ_io_enq_bits_addr; // @[VeriAXIRam.scala 34:22]
  wire [3:0] instRQ_io_enq_bits_len; // @[VeriAXIRam.scala 34:22]
  wire [1:0] instRQ_io_enq_bits_burst; // @[VeriAXIRam.scala 34:22]
  wire  instRQ_io_deq_ready; // @[VeriAXIRam.scala 34:22]
  wire  instRQ_io_deq_valid; // @[VeriAXIRam.scala 34:22]
  wire [31:0] instRQ_io_deq_bits_addr; // @[VeriAXIRam.scala 34:22]
  wire [3:0] instRQ_io_deq_bits_len; // @[VeriAXIRam.scala 34:22]
  wire [1:0] instRQ_io_deq_bits_burst; // @[VeriAXIRam.scala 34:22]
  wire  dataRQ_clock; // @[VeriAXIRam.scala 35:22]
  wire  dataRQ_reset; // @[VeriAXIRam.scala 35:22]
  wire  dataRQ_io_enq_ready; // @[VeriAXIRam.scala 35:22]
  wire  dataRQ_io_enq_valid; // @[VeriAXIRam.scala 35:22]
  wire [31:0] dataRQ_io_enq_bits_addr; // @[VeriAXIRam.scala 35:22]
  wire [3:0] dataRQ_io_enq_bits_len; // @[VeriAXIRam.scala 35:22]
  wire [1:0] dataRQ_io_enq_bits_burst; // @[VeriAXIRam.scala 35:22]
  wire  dataRQ_io_deq_ready; // @[VeriAXIRam.scala 35:22]
  wire  dataRQ_io_deq_valid; // @[VeriAXIRam.scala 35:22]
  wire [31:0] dataRQ_io_deq_bits_addr; // @[VeriAXIRam.scala 35:22]
  wire [3:0] dataRQ_io_deq_bits_len; // @[VeriAXIRam.scala 35:22]
  wire [1:0] dataRQ_io_deq_bits_burst; // @[VeriAXIRam.scala 35:22]
  wire  dataWQ_clock; // @[VeriAXIRam.scala 47:22]
  wire  dataWQ_reset; // @[VeriAXIRam.scala 47:22]
  wire  dataWQ_io_enq_ready; // @[VeriAXIRam.scala 47:22]
  wire  dataWQ_io_enq_valid; // @[VeriAXIRam.scala 47:22]
  wire [31:0] dataWQ_io_enq_bits_addr; // @[VeriAXIRam.scala 47:22]
  wire [3:0] dataWQ_io_enq_bits_len; // @[VeriAXIRam.scala 47:22]
  wire [1:0] dataWQ_io_enq_bits_burst; // @[VeriAXIRam.scala 47:22]
  wire  dataWQ_io_deq_ready; // @[VeriAXIRam.scala 47:22]
  wire  dataWQ_io_deq_valid; // @[VeriAXIRam.scala 47:22]
  wire [31:0] dataWQ_io_deq_bits_addr; // @[VeriAXIRam.scala 47:22]
  wire [3:0] dataWQ_io_deq_bits_len; // @[VeriAXIRam.scala 47:22]
  wire [1:0] dataWQ_io_deq_bits_burst; // @[VeriAXIRam.scala 47:22]
  reg  rState; // @[VeriAXIRam.scala 33:23]
  wire  currentID = instRQ_io_deq_valid ? 1'h0 : 1'h1; // @[VeriAXIRam.scala 36:22]
  reg [1:0] rBurst; // @[VeriAXIRam.scala 38:23]
  reg [3:0] rLen; // @[VeriAXIRam.scala 39:21]
  reg [2:0] rWrapSel; // @[VeriAXIRam.scala 40:25]
  reg [31:0] rRamAddr; // @[VeriAXIRam.scala 41:25]
  reg [1:0] wState; // @[VeriAXIRam.scala 46:23]
  wire  _T_36 = ~rState; // @[Conditional.scala 37:30]
  wire  _T_37 = 4'h1 == instRQ_io_deq_bits_len; // @[Mux.scala 80:60]
  wire [1:0] _T_38 = _T_37 ? 2'h3 : 2'h0; // @[Mux.scala 80:57]
  wire  _T_39 = 4'h3 == instRQ_io_deq_bits_len; // @[Mux.scala 80:60]
  wire  _T_41 = 4'h7 == instRQ_io_deq_bits_len; // @[Mux.scala 80:60]
  wire  _T_43 = 4'hf == instRQ_io_deq_bits_len; // @[Mux.scala 80:60]
  wire  _T_45 = 4'h1 == dataRQ_io_deq_bits_len; // @[Mux.scala 80:60]
  wire [1:0] _T_46 = _T_45 ? 2'h3 : 2'h0; // @[Mux.scala 80:57]
  wire  _T_47 = 4'h3 == dataRQ_io_deq_bits_len; // @[Mux.scala 80:60]
  wire  _T_49 = 4'h7 == dataRQ_io_deq_bits_len; // @[Mux.scala 80:60]
  wire  _T_51 = 4'hf == dataRQ_io_deq_bits_len; // @[Mux.scala 80:60]
  wire  _GEN_5 = dataRQ_io_deq_ready | rState; // @[VeriAXIRam.scala 55:39]
  wire  _GEN_11 = instRQ_io_deq_ready | _GEN_5; // @[VeriAXIRam.scala 51:33]
  wire  _T_54 = rLen == 4'h0; // @[VeriAXIRam.scala 63:19]
  wire [31:0] _T_56 = rRamAddr + 32'h4; // @[VeriAXIRam.scala 115:26]
  wire [31:0] _T_57 = rRamAddr >> rWrapSel; // @[VeriAXIRam.scala 117:57]
  wire [38:0] _GEN_54 = {{7'd0}, _T_57}; // @[VeriAXIRam.scala 117:70]
  wire [38:0] _T_58 = _GEN_54 << rWrapSel; // @[VeriAXIRam.scala 117:70]
  wire [5:0] _GEN_55 = {{3'd0}, rWrapSel}; // @[VeriAXIRam.scala 120:40]
  wire [5:0] _T_62 = 6'h20 - _GEN_55; // @[VeriAXIRam.scala 120:40]
  wire [94:0] _GEN_56 = {{63'd0}, _T_56}; // @[VeriAXIRam.scala 120:31]
  wire [94:0] _T_63 = _GEN_56 << _T_62; // @[VeriAXIRam.scala 120:31]
  wire [31:0] low = _T_63[31:0] >> _T_62; // @[VeriAXIRam.scala 120:69]
  wire [31:0] high = _T_58[31:0];
  wire [31:0] _T_68 = high | low; // @[VeriAXIRam.scala 122:16]
  wire  _T_69 = 2'h1 == rBurst; // @[Mux.scala 80:60]
  wire  _T_71 = 2'h2 == rBurst; // @[Mux.scala 80:60]
  wire [3:0] _T_74 = rLen - 4'h1; // @[VeriAXIRam.scala 67:24]
  wire  _T_79 = _T_36 & instRQ_io_deq_valid; // @[VeriAXIRam.scala 75:44]
  wire  _T_80 = ~currentID; // @[VeriAXIRam.scala 75:80]
  wire  _T_86 = _T_36 & dataRQ_io_deq_valid; // @[VeriAXIRam.scala 79:44]
  reg [31:0] wRamAddr; // @[VeriAXIRam.scala 90:25]
  wire  _T_95 = 2'h0 == wState; // @[Conditional.scala 37:30]
  wire [29:0] addr = wRamAddr[31:2]; // @[VeriAXIRam.scala 164:26]
  wire [15:0] _T_152 = {mem_internalData_data[15:8],mem_internalData_data[7:0]}; // @[Cat.scala 29:58]
  wire [15:0] _T_153 = {mem_internalData_data[31:24],mem_internalData_data[23:16]}; // @[Cat.scala 29:58]
  wire  _T_159 = wState == 2'h0; // @[VeriAXIRam.scala 173:33]
  Queue instRQ ( // @[VeriAXIRam.scala 34:22]
    .clock(instRQ_clock),
    .reset(instRQ_reset),
    .io_enq_ready(instRQ_io_enq_ready),
    .io_enq_valid(instRQ_io_enq_valid),
    .io_enq_bits_addr(instRQ_io_enq_bits_addr),
    .io_enq_bits_len(instRQ_io_enq_bits_len),
    .io_enq_bits_burst(instRQ_io_enq_bits_burst),
    .io_deq_ready(instRQ_io_deq_ready),
    .io_deq_valid(instRQ_io_deq_valid),
    .io_deq_bits_addr(instRQ_io_deq_bits_addr),
    .io_deq_bits_len(instRQ_io_deq_bits_len),
    .io_deq_bits_burst(instRQ_io_deq_bits_burst)
  );
  Queue dataRQ ( // @[VeriAXIRam.scala 35:22]
    .clock(dataRQ_clock),
    .reset(dataRQ_reset),
    .io_enq_ready(dataRQ_io_enq_ready),
    .io_enq_valid(dataRQ_io_enq_valid),
    .io_enq_bits_addr(dataRQ_io_enq_bits_addr),
    .io_enq_bits_len(dataRQ_io_enq_bits_len),
    .io_enq_bits_burst(dataRQ_io_enq_bits_burst),
    .io_deq_ready(dataRQ_io_deq_ready),
    .io_deq_valid(dataRQ_io_deq_valid),
    .io_deq_bits_addr(dataRQ_io_deq_bits_addr),
    .io_deq_bits_len(dataRQ_io_deq_bits_len),
    .io_deq_bits_burst(dataRQ_io_deq_bits_burst)
  );
  Queue dataWQ ( // @[VeriAXIRam.scala 47:22]
    .clock(dataWQ_clock),
    .reset(dataWQ_reset),
    .io_enq_ready(dataWQ_io_enq_ready),
    .io_enq_valid(dataWQ_io_enq_valid),
    .io_enq_bits_addr(dataWQ_io_enq_bits_addr),
    .io_enq_bits_len(dataWQ_io_enq_bits_len),
    .io_enq_bits_burst(dataWQ_io_enq_bits_burst),
    .io_deq_ready(dataWQ_io_deq_ready),
    .io_deq_valid(dataWQ_io_deq_valid),
    .io_deq_bits_addr(dataWQ_io_deq_bits_addr),
    .io_deq_bits_len(dataWQ_io_deq_bits_len),
    .io_deq_bits_burst(dataWQ_io_deq_bits_burst)
  );
  assign mem__T_92_addr = rRamAddr[13:2];
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign mem__T_92_data = mem[mem__T_92_addr]; // @[VeriAXIRam.scala 21:16]
  `else
  assign mem__T_92_data = mem__T_92_addr >= 12'hfff ? _RAND_1[31:0] : mem[mem__T_92_addr]; // @[VeriAXIRam.scala 21:16]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign mem_internalData_addr = addr[11:0];
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign mem_internalData_data = mem[mem_internalData_addr]; // @[VeriAXIRam.scala 21:16]
  `else
  assign mem_internalData_data = mem_internalData_addr >= 12'hfff ? _RAND_2[31:0] : mem[mem_internalData_addr]; // @[VeriAXIRam.scala 21:16]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign mem__T_155_data = {_T_153,_T_152};
  assign mem__T_155_addr = addr[11:0];
  assign mem__T_155_mask = 1'h1;
  assign mem__T_155_en = 1'h0;
  assign io_axi_ar_ready = instRQ_io_enq_ready & dataRQ_io_enq_ready; // @[VeriAXIRam.scala 81:12]
  assign io_axi_r_valid = rState; // @[VeriAXIRam.scala 86:11]
  assign io_axi_r_bits_data = mem__T_92_data; // @[VeriAXIRam.scala 83:15]
  assign io_axi_r_bits_last = rLen == 4'h0; // @[VeriAXIRam.scala 85:15]
  assign instRQ_clock = clock;
  assign instRQ_reset = reset;
  assign instRQ_io_enq_valid = io_axi_ar_ready & io_axi_ar_valid; // @[VeriAXIRam.scala 73:23]
  assign instRQ_io_enq_bits_addr = io_axi_ar_bits_addr; // @[VeriAXIRam.scala 74:22]
  assign instRQ_io_enq_bits_len = 4'h1; // @[VeriAXIRam.scala 74:22]
  assign instRQ_io_enq_bits_burst = 2'h2; // @[VeriAXIRam.scala 74:22]
  assign instRQ_io_deq_ready = _T_79 & _T_80; // @[VeriAXIRam.scala 75:23]
  assign dataRQ_clock = clock;
  assign dataRQ_reset = reset;
  assign dataRQ_io_enq_valid = 1'h0; // @[VeriAXIRam.scala 77:23]
  assign dataRQ_io_enq_bits_addr = io_axi_ar_bits_addr; // @[VeriAXIRam.scala 78:22]
  assign dataRQ_io_enq_bits_len = 4'h1; // @[VeriAXIRam.scala 78:22]
  assign dataRQ_io_enq_bits_burst = 2'h2; // @[VeriAXIRam.scala 78:22]
  assign dataRQ_io_deq_ready = _T_86 & currentID; // @[VeriAXIRam.scala 79:23]
  assign dataWQ_clock = clock;
  assign dataWQ_reset = reset;
  assign dataWQ_io_enq_valid = 1'h0; // @[VeriAXIRam.scala 171:23]
  assign dataWQ_io_enq_bits_addr = 32'h0; // @[VeriAXIRam.scala 172:22]
  assign dataWQ_io_enq_bits_len = 4'h0; // @[VeriAXIRam.scala 172:22]
  assign dataWQ_io_enq_bits_burst = 2'h0; // @[VeriAXIRam.scala 172:22]
  assign dataWQ_io_deq_ready = _T_159 & dataWQ_io_deq_valid; // @[VeriAXIRam.scala 173:23]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_GARBAGE_ASSIGN
  _RAND_1 = {1{`RANDOM}};
  _RAND_2 = {1{`RANDOM}};
`endif // RANDOMIZE_GARBAGE_ASSIGN
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4095; initvar = initvar+1)
    mem[initvar] = _RAND_0[31:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  rState = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  rBurst = _RAND_4[1:0];
  _RAND_5 = {1{`RANDOM}};
  rLen = _RAND_5[3:0];
  _RAND_6 = {1{`RANDOM}};
  rWrapSel = _RAND_6[2:0];
  _RAND_7 = {1{`RANDOM}};
  rRamAddr = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  wState = _RAND_8[1:0];
  _RAND_9 = {1{`RANDOM}};
  wRamAddr = _RAND_9[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(mem__T_155_en & mem__T_155_mask) begin
      mem[mem__T_155_addr] <= mem__T_155_data; // @[VeriAXIRam.scala 21:16]
    end
    if (reset) begin
      rState <= 1'h0;
    end else if (_T_36) begin
      rState <= _GEN_11;
    end else if (rState) begin
      if (io_axi_r_ready) begin
        if (_T_54) begin
          rState <= 1'h0;
        end
      end
    end
    if (reset) begin
      rBurst <= 2'h0;
    end else if (_T_36) begin
      if (instRQ_io_deq_ready) begin
        rBurst <= instRQ_io_deq_bits_burst;
      end else if (dataRQ_io_deq_ready) begin
        rBurst <= dataRQ_io_deq_bits_burst;
      end
    end
    if (reset) begin
      rLen <= 4'h0;
    end else if (_T_36) begin
      if (instRQ_io_deq_ready) begin
        rLen <= instRQ_io_deq_bits_len;
      end else if (dataRQ_io_deq_ready) begin
        rLen <= dataRQ_io_deq_bits_len;
      end
    end else if (rState) begin
      if (io_axi_r_ready) begin
        if (!(_T_54)) begin
          rLen <= _T_74;
        end
      end
    end
    if (reset) begin
      rWrapSel <= 3'h0;
    end else if (_T_36) begin
      if (instRQ_io_deq_ready) begin
        if (_T_43) begin
          rWrapSel <= 3'h6;
        end else if (_T_41) begin
          rWrapSel <= 3'h5;
        end else if (_T_39) begin
          rWrapSel <= 3'h4;
        end else begin
          rWrapSel <= {{1'd0}, _T_38};
        end
      end else if (dataRQ_io_deq_ready) begin
        if (_T_51) begin
          rWrapSel <= 3'h6;
        end else if (_T_49) begin
          rWrapSel <= 3'h5;
        end else if (_T_47) begin
          rWrapSel <= 3'h4;
        end else begin
          rWrapSel <= {{1'd0}, _T_46};
        end
      end
    end
    if (reset) begin
      rRamAddr <= 32'h0;
    end else if (_T_36) begin
      if (instRQ_io_deq_ready) begin
        rRamAddr <= instRQ_io_deq_bits_addr;
      end else if (dataRQ_io_deq_ready) begin
        rRamAddr <= dataRQ_io_deq_bits_addr;
      end
    end else if (rState) begin
      if (io_axi_r_ready) begin
        if (!(_T_54)) begin
          if (_T_71) begin
            rRamAddr <= _T_68;
          end else if (_T_69) begin
            rRamAddr <= _T_56;
          end else begin
            rRamAddr <= 32'h0;
          end
        end
      end
    end
    if (reset) begin
      wState <= 2'h0;
    end else if (_T_95) begin
      if (dataWQ_io_deq_valid) begin
        wState <= 2'h1;
      end
    end
    if (reset) begin
      wRamAddr <= 32'h0;
    end else if (_T_95) begin
      if (dataWQ_io_deq_valid) begin
        wRamAddr <= dataWQ_io_deq_bits_addr;
      end
    end
  end
endmodule
module ICacheVeri(
  input         clock,
  input         reset,
  output        io_addr_ready,
  input         io_addr_valid,
  input  [31:0] io_addr_bits,
  input         io_data_ready,
  output        io_data_valid,
  output [31:0] io_data_bits,
  input         io_flush
);
  wire  insCache_clock; // @[InstrCache.scala 109:26]
  wire  insCache_reset; // @[InstrCache.scala 109:26]
  wire  insCache_io_addr_ready; // @[InstrCache.scala 109:26]
  wire  insCache_io_addr_valid; // @[InstrCache.scala 109:26]
  wire [31:0] insCache_io_addr_bits; // @[InstrCache.scala 109:26]
  wire  insCache_io_data_ready; // @[InstrCache.scala 109:26]
  wire  insCache_io_data_valid; // @[InstrCache.scala 109:26]
  wire [31:0] insCache_io_data_bits; // @[InstrCache.scala 109:26]
  wire  insCache_io_flush; // @[InstrCache.scala 109:26]
  wire  insCache_io_axi_ar_ready; // @[InstrCache.scala 109:26]
  wire  insCache_io_axi_ar_valid; // @[InstrCache.scala 109:26]
  wire [31:0] insCache_io_axi_ar_bits_addr; // @[InstrCache.scala 109:26]
  wire  insCache_io_axi_r_ready; // @[InstrCache.scala 109:26]
  wire  insCache_io_axi_r_valid; // @[InstrCache.scala 109:26]
  wire [31:0] insCache_io_axi_r_bits_data; // @[InstrCache.scala 109:26]
  wire  insCache_io_axi_r_bits_last; // @[InstrCache.scala 109:26]
  wire  ram_clock; // @[InstrCache.scala 110:26]
  wire  ram_reset; // @[InstrCache.scala 110:26]
  wire  ram_io_axi_ar_ready; // @[InstrCache.scala 110:26]
  wire  ram_io_axi_ar_valid; // @[InstrCache.scala 110:26]
  wire [31:0] ram_io_axi_ar_bits_addr; // @[InstrCache.scala 110:26]
  wire  ram_io_axi_r_ready; // @[InstrCache.scala 110:26]
  wire  ram_io_axi_r_valid; // @[InstrCache.scala 110:26]
  wire [31:0] ram_io_axi_r_bits_data; // @[InstrCache.scala 110:26]
  wire  ram_io_axi_r_bits_last; // @[InstrCache.scala 110:26]
  InstrCache insCache ( // @[InstrCache.scala 109:26]
    .clock(insCache_clock),
    .reset(insCache_reset),
    .io_addr_ready(insCache_io_addr_ready),
    .io_addr_valid(insCache_io_addr_valid),
    .io_addr_bits(insCache_io_addr_bits),
    .io_data_ready(insCache_io_data_ready),
    .io_data_valid(insCache_io_data_valid),
    .io_data_bits(insCache_io_data_bits),
    .io_flush(insCache_io_flush),
    .io_axi_ar_ready(insCache_io_axi_ar_ready),
    .io_axi_ar_valid(insCache_io_axi_ar_valid),
    .io_axi_ar_bits_addr(insCache_io_axi_ar_bits_addr),
    .io_axi_r_ready(insCache_io_axi_r_ready),
    .io_axi_r_valid(insCache_io_axi_r_valid),
    .io_axi_r_bits_data(insCache_io_axi_r_bits_data),
    .io_axi_r_bits_last(insCache_io_axi_r_bits_last)
  );
  VeriAXIRam ram ( // @[InstrCache.scala 110:26]
    .clock(ram_clock),
    .reset(ram_reset),
    .io_axi_ar_ready(ram_io_axi_ar_ready),
    .io_axi_ar_valid(ram_io_axi_ar_valid),
    .io_axi_ar_bits_addr(ram_io_axi_ar_bits_addr),
    .io_axi_r_ready(ram_io_axi_r_ready),
    .io_axi_r_valid(ram_io_axi_r_valid),
    .io_axi_r_bits_data(ram_io_axi_r_bits_data),
    .io_axi_r_bits_last(ram_io_axi_r_bits_last)
  );
  assign io_addr_ready = insCache_io_addr_ready; // @[InstrCache.scala 112:39]
  assign io_data_valid = insCache_io_data_valid; // @[InstrCache.scala 113:39]
  assign io_data_bits = insCache_io_data_bits; // @[InstrCache.scala 113:39]
  assign insCache_clock = clock;
  assign insCache_reset = reset;
  assign insCache_io_addr_valid = io_addr_valid; // @[InstrCache.scala 112:39]
  assign insCache_io_addr_bits = io_addr_bits; // @[InstrCache.scala 112:39]
  assign insCache_io_data_ready = io_data_ready; // @[InstrCache.scala 113:39]
  assign insCache_io_flush = io_flush; // @[InstrCache.scala 114:39]
  assign insCache_io_axi_ar_ready = ram_io_axi_ar_ready; // @[InstrCache.scala 111:39]
  assign insCache_io_axi_r_valid = ram_io_axi_r_valid; // @[InstrCache.scala 111:39]
  assign insCache_io_axi_r_bits_data = ram_io_axi_r_bits_data; // @[InstrCache.scala 111:39]
  assign insCache_io_axi_r_bits_last = ram_io_axi_r_bits_last; // @[InstrCache.scala 111:39]
  assign ram_clock = clock;
  assign ram_reset = reset;
  assign ram_io_axi_ar_valid = insCache_io_axi_ar_valid; // @[InstrCache.scala 111:39]
  assign ram_io_axi_ar_bits_addr = insCache_io_axi_ar_bits_addr; // @[InstrCache.scala 111:39]
  assign ram_io_axi_r_ready = insCache_io_axi_r_ready; // @[InstrCache.scala 111:39]
endmodule
